<?xml version="1.0" encoding="utf-8" ?>
<svg baseProfile="full" height="1500" version="1.1" width="1500" xmlns="http://www.w3.org/2000/svg" xmlns:ev="http://www.w3.org/2001/xml-events" xmlns:xlink="http://www.w3.org/1999/xlink"><defs><linearGradient id="ropegrad" x1="0%" x2="100%" y1="0%" y2="100%"><stop offset="0" stop-color="#000000" /><stop offset="1" stop-color="#000000" /></linearGradient><filter height="140%" id="glow" width="140%" x="-20%" y="-20%"><feGaussianBlur in="SourceGraphic" result="blur" stdDeviation="2" /><feColorMatrix in="blur" result="soft" type="matrix" values="[0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9, 0]" /><feMerge><feMergeNode in="soft" /><feMergeNode in="SourceGraphic" /></feMerge></filter><filter height="140%" id="emboss" width="140%" x="-20%" y="-20%"><feGaussianBlur in="SourceAlpha" result="alpha" stdDeviation="0.7" /><feSpecularLighting in="alpha" lighting-color="#ffffff" result="spec" specularConstant="0.6" specularExponent="15" surfaceScale="2"><fePointLight x="0" y="-5000" z="2000" /></feSpecularLighting><feComposite in="spec" in2="SourceGraphic" operator="in" result="lit" /><feMerge><feMergeNode in="lit" /><feMergeNode in="SourceGraphic" /></feMerge></filter><filter height="100%" id="paper" width="100%" x="0%" y="0%"><feTurbulence baseFrequency="0.8" numOctaves="2" result="noise" seed="3" type="fractalNoise" /><feColorMatrix in="noise" result="grain" type="saturate" values="0.15" /><feBlend in="SourceGraphic" in2="grain" mode="multiply" /></filter><radialGradient cx="50%" cy="50%" id="vign" r="65%"><stop offset="0" stop-color="#ffffff" /><stop offset="1" stop-color="#ffffff" /></radialGradient></defs><g><rect fill="#ffffff" height="1500" width="1500" x="0" y="0" /><rect fill="url(#vign)" filter="url(#paper)" height="1500" width="1500" x="0" y="0" /></g><g><rect fill="none" height="1496" stroke="#000000" stroke-width="4" width="1496" x="2" y="2" /><circle cx="72.0" cy="72.0" fill="#000000" opacity="0.9" r="26.4" /><g><path d="M 72.00,72.00 Q 81.81,77.66 92.59,72.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 79.28,80.68 91.35,79.04" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 75.87,82.64 87.77,85.24" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 72.00,83.33 82.30,89.83" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 68.13,82.64 75.58,92.28" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 64.72,80.68 68.42,92.28" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 62.19,77.66 61.70,89.83" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 60.85,73.97 56.23,85.24" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 60.85,70.03 52.65,79.04" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 62.19,66.34 51.41,72.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 64.72,63.32 52.65,64.96" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 68.13,61.36 56.23,58.76" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 72.00,60.67 61.70,54.17" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 75.87,61.36 68.42,51.72" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 79.28,63.32 75.58,51.72" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 81.81,66.34 82.30,54.17" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 83.15,70.03 87.77,58.76" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,72.00 Q 83.15,73.97 91.35,64.96" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /></g><circle cx="1428.0" cy="72.0" fill="#000000" opacity="0.9" r="26.4" /><g><path d="M 1428.00,72.00 Q 1437.81,77.66 1448.59,72.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1435.28,80.68 1447.35,79.04" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1431.87,82.64 1443.77,85.24" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1428.00,83.33 1438.30,89.83" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1424.13,82.64 1431.58,92.28" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1420.72,80.68 1424.42,92.28" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1418.19,77.66 1417.70,89.83" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1416.85,73.97 1412.23,85.24" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1416.85,70.03 1408.65,79.04" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1418.19,66.34 1407.41,72.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1420.72,63.32 1408.65,64.96" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1424.13,61.36 1412.23,58.76" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1428.00,60.67 1417.70,54.17" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1431.87,61.36 1424.42,51.72" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1435.28,63.32 1431.58,51.72" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1437.81,66.34 1438.30,54.17" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1439.15,70.03 1443.77,58.76" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 1428.00,72.00 Q 1439.15,73.97 1447.35,64.96" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /></g><circle cx="72.0" cy="1428.0" fill="#000000" opacity="0.9" r="26.4" /><g><path d="M 72.00,1428.00 Q 81.81,1433.66 92.59,1428.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 79.28,1436.68 91.35,1435.04" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 75.87,1438.64 87.77,1441.24" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 72.00,1439.33 82.30,1445.83" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 68.13,1438.64 75.58,1448.28" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 64.72,1436.68 68.42,1448.28" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 62.19,1433.66 61.70,1445.83" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 60.85,1429.97 56.23,1441.24" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 60.85,1426.03 52.65,1435.04" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 62.19,1422.34 51.41,1428.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 64.72,1419.32 52.65,1420.96" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 68.13,1417.36 56.23,1414.76" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 72.00,1416.67 61.70,1410.17" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 75.87,1417.36 68.42,1407.72" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 79.28,1419.32 75.58,1407.72" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 81.81,1422.34 82.30,1410.17" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 83.15,1426.03 87.77,1414.76" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /><path d="M 72.00,1428.00 Q 83.15,1429.97 91.35,1420.96" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="1.2" /></g><g opacity="0.3"><circle cx="120.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="120.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="120.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="144.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="144.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="168.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="168.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="192.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="192.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="216.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="216.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="240.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="240.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="264.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="264.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="288.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="288.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="312.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="312.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="336.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="336.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="360.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="360.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="384.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="384.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="408.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="408.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="432.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="432.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="456.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="456.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="480.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="480.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="504.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="504.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="528.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="528.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="552.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="552.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="576.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="576.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="600.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="600.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="624.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="624.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="648.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="648.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="672.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="672.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="696.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="696.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="720.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="720.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="744.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="744.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="768.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="768.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="792.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="792.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="816.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="816.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="840.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="840.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="864.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="864.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="888.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="888.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="912.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="912.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="936.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="936.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="960.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="960.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="984.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="984.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1008.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1008.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1032.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1032.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1056.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1056.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1080.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1080.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1104.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1104.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1128.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1128.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1152.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1152.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1176.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1176.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1200.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1200.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1224.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1224.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1248.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1248.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1272.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1272.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1296.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1296.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1320.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1320.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1344.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1344.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="120.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="120.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="144.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="144.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="168.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="168.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="192.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="192.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="216.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="216.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="240.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="240.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="264.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="264.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="288.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="288.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="312.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="312.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="336.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="336.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="360.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="360.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="384.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="384.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="408.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="408.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="432.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="432.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="456.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="456.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="480.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="480.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="504.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="504.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="528.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="528.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="552.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="552.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="576.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="576.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="600.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="600.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="624.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="624.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="648.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="648.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="672.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="672.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="696.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="696.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="720.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="720.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="744.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="744.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="768.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="768.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="792.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="792.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="816.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="816.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="840.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="840.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="864.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="864.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="888.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="888.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="912.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="912.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="936.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="936.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="960.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="960.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="984.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="984.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1008.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1008.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1032.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1032.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1056.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1056.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1080.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1080.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1104.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1104.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1128.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1128.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1152.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1152.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1176.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1176.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1200.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1200.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1224.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1224.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1248.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1248.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1272.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1272.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1296.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1296.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1320.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1320.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1344.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1344.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /><circle cx="1368.0" cy="1368.0" fill="#666666" opacity="0.9" r="5.4" /><circle cx="1368.0" cy="1368.0" fill="none" opacity="0.6" r="3.5999999999999996" stroke="#666666" stroke-width="0.5" /></g></g><g><path d="M 124.80,150.00 C 135.78,139.02 146.58,128.22 150.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 175.20,150.00 C 164.22,160.98 153.42,171.78 150.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 150.00,134.88 C 156.40,141.28 163.26,148.14 165.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,165.12 C 143.60,158.72 136.74,151.86 134.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 184.80,150.00 C 195.78,139.02 206.58,128.22 210.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 235.20,150.00 C 224.22,160.98 213.42,171.78 210.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,134.88 C 216.40,141.28 223.26,148.14 225.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,165.12 C 203.60,158.72 196.74,151.86 194.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,124.80 C 280.98,135.78 291.78,146.58 295.20,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,175.20 C 259.02,164.22 248.22,153.42 244.80,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 285.12,150.00 C 278.72,156.40 271.86,163.26 270.00,165.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 254.88,150.00 C 261.28,143.60 268.14,136.74 270.00,134.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,150.00 C 315.78,139.02 326.58,128.22 330.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,150.00 C 344.22,160.98 333.42,171.78 330.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 330.00,134.88 C 336.40,141.28 343.26,148.14 345.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,165.12 C 323.60,158.72 316.74,151.86 314.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,150.00 C 375.78,139.02 386.58,128.22 390.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,150.00 C 404.22,160.98 393.42,171.78 390.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 390.00,134.88 C 396.40,141.28 403.26,148.14 405.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,165.12 C 383.60,158.72 376.74,151.86 374.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 450.00,175.20 C 439.02,164.22 428.22,153.42 424.80,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,124.80 C 460.98,135.78 471.78,146.58 475.20,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 434.88,150.00 C 441.28,143.60 448.14,136.74 450.00,134.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 465.12,150.00 C 458.72,156.40 451.86,163.26 450.00,165.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,175.20 C 499.02,164.22 488.22,153.42 484.80,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,124.80 C 520.98,135.78 531.78,146.58 535.20,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,150.00 Q 517.32,153.03 523.20,150.00 Q 517.32,146.97 510.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,150.00 Q 513.03,157.32 519.33,159.33 Q 517.32,153.03 510.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,150.00 Q 506.97,157.32 510.00,163.20 Q 513.03,157.32 510.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,150.00 Q 502.68,153.03 500.67,159.33 Q 506.97,157.32 510.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,150.00 Q 502.68,146.97 496.80,150.00 Q 502.68,153.03 510.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,150.00 Q 506.97,142.68 500.67,140.67 Q 502.68,146.97 510.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,150.00 Q 513.03,142.68 510.00,136.80 Q 506.97,142.68 510.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,150.00 Q 517.32,146.97 519.33,140.67 Q 513.03,142.68 510.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,150.00 Q 510.93,153.48 515.09,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,150.00 Q 506.52,150.93 504.91,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,150.00 Q 509.07,146.52 504.91,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,150.00 Q 513.48,149.07 515.09,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="150.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 494.88,150.00 C 501.28,143.60 508.14,136.74 510.00,134.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 525.12,150.00 C 518.72,156.40 511.86,163.26 510.00,165.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,150.00 C 555.78,139.02 566.58,128.22 570.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,150.00 C 584.22,160.98 573.42,171.78 570.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 570.00,150.00 Q 577.32,153.03 583.20,150.00 Q 577.32,146.97 570.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,150.00 Q 573.03,157.32 579.33,159.33 Q 577.32,153.03 570.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,150.00 Q 566.97,157.32 570.00,163.20 Q 573.03,157.32 570.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,150.00 Q 562.68,153.03 560.67,159.33 Q 566.97,157.32 570.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,150.00 Q 562.68,146.97 556.80,150.00 Q 562.68,153.03 570.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,150.00 Q 566.97,142.68 560.67,140.67 Q 562.68,146.97 570.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,150.00 Q 573.03,142.68 570.00,136.80 Q 566.97,142.68 570.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,150.00 Q 577.32,146.97 579.33,140.67 Q 573.03,142.68 570.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,150.00 Q 570.93,153.48 575.09,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,150.00 Q 566.52,150.93 564.91,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,150.00 Q 569.07,146.52 564.91,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,150.00 Q 573.48,149.07 575.09,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="570.0" cy="150.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 570.00,134.88 C 576.40,141.28 583.26,148.14 585.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,165.12 C 563.60,158.72 556.74,151.86 554.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,150.00 C 615.78,139.02 626.58,128.22 630.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,150.00 C 644.22,160.98 633.42,171.78 630.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,134.88 C 636.40,141.28 643.26,148.14 645.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,165.12 C 623.60,158.72 616.74,151.86 614.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 664.80,150.00 C 675.78,139.02 686.58,128.22 690.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 715.20,150.00 C 704.22,160.98 693.42,171.78 690.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 690.00,134.88 C 696.40,141.28 703.26,148.14 705.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,165.12 C 683.60,158.72 676.74,151.86 674.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 724.80,150.00 C 735.78,139.02 746.58,128.22 750.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 775.20,150.00 C 764.22,160.98 753.42,171.78 750.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,134.88 C 756.40,141.28 763.26,148.14 765.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,165.12 C 743.60,158.72 736.74,151.86 734.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 784.80,150.00 C 795.78,139.02 806.58,128.22 810.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 835.20,150.00 C 824.22,160.98 813.42,171.78 810.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,134.88 C 816.40,141.28 823.26,148.14 825.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,165.12 C 803.60,158.72 796.74,151.86 794.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 844.80,150.00 C 855.78,139.02 866.58,128.22 870.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 895.20,150.00 C 884.22,160.98 873.42,171.78 870.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 870.00,134.88 C 876.40,141.28 883.26,148.14 885.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,165.12 C 863.60,158.72 856.74,151.86 854.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 904.80,150.00 C 915.78,139.02 926.58,128.22 930.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 955.20,150.00 C 944.22,160.98 933.42,171.78 930.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 930.00,134.88 C 936.40,141.28 943.26,148.14 945.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,165.12 C 923.60,158.72 916.74,151.86 914.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 964.80,150.00 C 975.78,139.02 986.58,128.22 990.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1015.20,150.00 C 1004.22,160.98 993.42,171.78 990.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 990.00,134.88 C 996.40,141.28 1003.26,148.14 1005.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,165.12 C 983.60,158.72 976.74,151.86 974.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,150.00 C 1035.78,139.02 1046.58,128.22 1050.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,150.00 C 1064.22,160.98 1053.42,171.78 1050.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,134.88 C 1056.40,141.28 1063.26,148.14 1065.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,165.12 C 1043.60,158.72 1036.74,151.86 1034.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1110.00,124.80 C 1120.98,135.78 1131.78,146.58 1135.20,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,175.20 C 1099.02,164.22 1088.22,153.42 1084.80,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1110.00,150.00 Q 1117.32,153.03 1123.20,150.00 Q 1117.32,146.97 1110.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,150.00 Q 1113.03,157.32 1119.33,159.33 Q 1117.32,153.03 1110.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,150.00 Q 1106.97,157.32 1110.00,163.20 Q 1113.03,157.32 1110.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,150.00 Q 1102.68,153.03 1100.67,159.33 Q 1106.97,157.32 1110.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,150.00 Q 1102.68,146.97 1096.80,150.00 Q 1102.68,153.03 1110.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,150.00 Q 1106.97,142.68 1100.67,140.67 Q 1102.68,146.97 1110.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,150.00 Q 1113.03,142.68 1110.00,136.80 Q 1106.97,142.68 1110.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,150.00 Q 1117.32,146.97 1119.33,140.67 Q 1113.03,142.68 1110.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,150.00 Q 1110.93,153.48 1115.09,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,150.00 Q 1106.52,150.93 1104.91,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,150.00 Q 1109.07,146.52 1104.91,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,150.00 Q 1113.48,149.07 1115.09,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1110.0" cy="150.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1125.12,150.00 C 1118.72,156.40 1111.86,163.26 1110.00,165.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1094.88,150.00 C 1101.28,143.60 1108.14,136.74 1110.00,134.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1170.00,175.20 C 1159.02,164.22 1148.22,153.42 1144.80,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,124.80 C 1180.98,135.78 1191.78,146.58 1195.20,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1154.88,150.00 C 1161.28,143.60 1168.14,136.74 1170.00,134.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1185.12,150.00 C 1178.72,156.40 1171.86,163.26 1170.00,165.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,175.20 C 1219.02,164.22 1208.22,153.42 1204.80,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,124.80 C 1240.98,135.78 1251.78,146.58 1255.20,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1214.88,150.00 C 1221.28,143.60 1228.14,136.74 1230.00,134.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1245.12,150.00 C 1238.72,156.40 1231.86,163.26 1230.00,165.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1315.20,150.00 C 1304.22,160.98 1293.42,171.78 1290.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1264.80,150.00 C 1275.78,139.02 1286.58,128.22 1290.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1290.00,150.00 Q 1297.32,153.03 1303.20,150.00 Q 1297.32,146.97 1290.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,150.00 Q 1293.03,157.32 1299.33,159.33 Q 1297.32,153.03 1290.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,150.00 Q 1286.97,157.32 1290.00,163.20 Q 1293.03,157.32 1290.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,150.00 Q 1282.68,153.03 1280.67,159.33 Q 1286.97,157.32 1290.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,150.00 Q 1282.68,146.97 1276.80,150.00 Q 1282.68,153.03 1290.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,150.00 Q 1286.97,142.68 1280.67,140.67 Q 1282.68,146.97 1290.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,150.00 Q 1293.03,142.68 1290.00,136.80 Q 1286.97,142.68 1290.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,150.00 Q 1297.32,146.97 1299.33,140.67 Q 1293.03,142.68 1290.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,150.00 Q 1290.93,153.48 1295.09,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,150.00 Q 1286.52,150.93 1284.91,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,150.00 Q 1289.07,146.52 1284.91,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,150.00 Q 1293.48,149.07 1295.09,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1290.0" cy="150.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1290.00,165.12 C 1283.60,158.72 1276.74,151.86 1274.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,134.88 C 1296.40,141.28 1303.26,148.14 1305.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1324.80,150.00 C 1335.78,139.02 1346.58,128.22 1350.00,124.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1375.20,150.00 C 1364.22,160.98 1353.42,171.78 1350.00,175.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1350.00,150.00 Q 1357.32,153.03 1363.20,150.00 Q 1357.32,146.97 1350.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,150.00 Q 1353.03,157.32 1359.33,159.33 Q 1357.32,153.03 1350.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,150.00 Q 1346.97,157.32 1350.00,163.20 Q 1353.03,157.32 1350.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,150.00 Q 1342.68,153.03 1340.67,159.33 Q 1346.97,157.32 1350.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,150.00 Q 1342.68,146.97 1336.80,150.00 Q 1342.68,153.03 1350.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,150.00 Q 1346.97,142.68 1340.67,140.67 Q 1342.68,146.97 1350.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,150.00 Q 1353.03,142.68 1350.00,136.80 Q 1346.97,142.68 1350.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,150.00 Q 1357.32,146.97 1359.33,140.67 Q 1353.03,142.68 1350.00,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,150.00 Q 1350.93,153.48 1355.09,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,150.00 Q 1346.52,150.93 1344.91,155.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,150.00 Q 1349.07,146.52 1344.91,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,150.00 Q 1353.48,149.07 1355.09,144.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1350.0" cy="150.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1350.00,134.88 C 1356.40,141.28 1363.26,148.14 1365.12,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,165.12 C 1343.60,158.72 1336.74,151.86 1334.88,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 175.20,210.00 C 164.22,220.98 153.42,231.78 150.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 124.80,210.00 C 135.78,199.02 146.58,188.22 150.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,210.00 Q 157.32,213.03 163.20,210.00 Q 157.32,206.97 150.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,210.00 Q 153.03,217.32 159.33,219.33 Q 157.32,213.03 150.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,210.00 Q 146.97,217.32 150.00,223.20 Q 153.03,217.32 150.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,210.00 Q 142.68,213.03 140.67,219.33 Q 146.97,217.32 150.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,210.00 Q 142.68,206.97 136.80,210.00 Q 142.68,213.03 150.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,210.00 Q 146.97,202.68 140.67,200.67 Q 142.68,206.97 150.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,210.00 Q 153.03,202.68 150.00,196.80 Q 146.97,202.68 150.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,210.00 Q 157.32,206.97 159.33,200.67 Q 153.03,202.68 150.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,210.00 Q 150.93,213.48 155.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,210.00 Q 146.52,210.93 144.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,210.00 Q 149.07,206.52 144.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,210.00 Q 153.48,209.07 155.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 150.00,225.12 C 143.60,218.72 136.74,211.86 134.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,194.88 C 156.40,201.28 163.26,208.14 165.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 210.00,235.20 C 199.02,224.22 188.22,213.42 184.80,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,184.80 C 220.98,195.78 231.78,206.58 235.20,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 194.88,210.00 C 201.28,203.60 208.14,196.74 210.00,194.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 225.12,210.00 C 218.72,216.40 211.86,223.26 210.00,225.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 295.20,210.00 C 284.22,220.98 273.42,231.78 270.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 244.80,210.00 C 255.78,199.02 266.58,188.22 270.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 270.00,210.00 Q 277.32,213.03 283.20,210.00 Q 277.32,206.97 270.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,210.00 Q 273.03,217.32 279.33,219.33 Q 277.32,213.03 270.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,210.00 Q 266.97,217.32 270.00,223.20 Q 273.03,217.32 270.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,210.00 Q 262.68,213.03 260.67,219.33 Q 266.97,217.32 270.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,210.00 Q 262.68,206.97 256.80,210.00 Q 262.68,213.03 270.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,210.00 Q 266.97,202.68 260.67,200.67 Q 262.68,206.97 270.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,210.00 Q 273.03,202.68 270.00,196.80 Q 266.97,202.68 270.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,210.00 Q 277.32,206.97 279.33,200.67 Q 273.03,202.68 270.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,210.00 Q 270.93,213.48 275.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,210.00 Q 266.52,210.93 264.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,210.00 Q 269.07,206.52 264.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,210.00 Q 273.48,209.07 275.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="270.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 270.00,225.12 C 263.60,218.72 256.74,211.86 254.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,194.88 C 276.40,201.28 283.26,208.14 285.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 330.00,184.80 C 340.98,195.78 351.78,206.58 355.20,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,235.20 C 319.02,224.22 308.22,213.42 304.80,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 330.00,210.00 Q 337.32,213.03 343.20,210.00 Q 337.32,206.97 330.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,210.00 Q 333.03,217.32 339.33,219.33 Q 337.32,213.03 330.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,210.00 Q 326.97,217.32 330.00,223.20 Q 333.03,217.32 330.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,210.00 Q 322.68,213.03 320.67,219.33 Q 326.97,217.32 330.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,210.00 Q 322.68,206.97 316.80,210.00 Q 322.68,213.03 330.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,210.00 Q 326.97,202.68 320.67,200.67 Q 322.68,206.97 330.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,210.00 Q 333.03,202.68 330.00,196.80 Q 326.97,202.68 330.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,210.00 Q 337.32,206.97 339.33,200.67 Q 333.03,202.68 330.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,210.00 Q 330.93,213.48 335.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,210.00 Q 326.52,210.93 324.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,210.00 Q 329.07,206.52 324.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,210.00 Q 333.48,209.07 335.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="330.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 345.12,210.00 C 338.72,216.40 331.86,223.26 330.00,225.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 314.88,210.00 C 321.28,203.60 328.14,196.74 330.00,194.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,210.00 C 375.78,199.02 386.58,188.22 390.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,210.00 C 404.22,220.98 393.42,231.78 390.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 390.00,194.88 C 396.40,201.28 403.26,208.14 405.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,225.12 C 383.60,218.72 376.74,211.86 374.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 475.20,210.00 C 464.22,220.98 453.42,231.78 450.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 424.80,210.00 C 435.78,199.02 446.58,188.22 450.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 450.00,225.12 C 443.60,218.72 436.74,211.86 434.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,194.88 C 456.40,201.28 463.26,208.14 465.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,235.20 C 499.02,224.22 488.22,213.42 484.80,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,184.80 C 520.98,195.78 531.78,206.58 535.20,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,210.00 Q 517.32,213.03 523.20,210.00 Q 517.32,206.97 510.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,210.00 Q 513.03,217.32 519.33,219.33 Q 517.32,213.03 510.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,210.00 Q 506.97,217.32 510.00,223.20 Q 513.03,217.32 510.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,210.00 Q 502.68,213.03 500.67,219.33 Q 506.97,217.32 510.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,210.00 Q 502.68,206.97 496.80,210.00 Q 502.68,213.03 510.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,210.00 Q 506.97,202.68 500.67,200.67 Q 502.68,206.97 510.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,210.00 Q 513.03,202.68 510.00,196.80 Q 506.97,202.68 510.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,210.00 Q 517.32,206.97 519.33,200.67 Q 513.03,202.68 510.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,210.00 Q 510.93,213.48 515.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,210.00 Q 506.52,210.93 504.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,210.00 Q 509.07,206.52 504.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,210.00 Q 513.48,209.07 515.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 494.88,210.00 C 501.28,203.60 508.14,196.74 510.00,194.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 525.12,210.00 C 518.72,216.40 511.86,223.26 510.00,225.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 570.00,184.80 C 580.98,195.78 591.78,206.58 595.20,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,235.20 C 559.02,224.22 548.22,213.42 544.80,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 585.12,210.00 C 578.72,216.40 571.86,223.26 570.00,225.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 554.88,210.00 C 561.28,203.60 568.14,196.74 570.00,194.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,210.00 C 615.78,199.02 626.58,188.22 630.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,210.00 C 644.22,220.98 633.42,231.78 630.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 630.00,210.00 Q 637.32,213.03 643.20,210.00 Q 637.32,206.97 630.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,210.00 Q 633.03,217.32 639.33,219.33 Q 637.32,213.03 630.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,210.00 Q 626.97,217.32 630.00,223.20 Q 633.03,217.32 630.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,210.00 Q 622.68,213.03 620.67,219.33 Q 626.97,217.32 630.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,210.00 Q 622.68,206.97 616.80,210.00 Q 622.68,213.03 630.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,210.00 Q 626.97,202.68 620.67,200.67 Q 622.68,206.97 630.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,210.00 Q 633.03,202.68 630.00,196.80 Q 626.97,202.68 630.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,210.00 Q 637.32,206.97 639.33,200.67 Q 633.03,202.68 630.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,210.00 Q 630.93,213.48 635.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,210.00 Q 626.52,210.93 624.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,210.00 Q 629.07,206.52 624.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,210.00 Q 633.48,209.07 635.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="630.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 630.00,194.88 C 636.40,201.28 643.26,208.14 645.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,225.12 C 623.60,218.72 616.74,211.86 614.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 715.20,210.00 C 704.22,220.98 693.42,231.78 690.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 664.80,210.00 C 675.78,199.02 686.58,188.22 690.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 690.00,210.00 Q 697.32,213.03 703.20,210.00 Q 697.32,206.97 690.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,210.00 Q 693.03,217.32 699.33,219.33 Q 697.32,213.03 690.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,210.00 Q 686.97,217.32 690.00,223.20 Q 693.03,217.32 690.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,210.00 Q 682.68,213.03 680.67,219.33 Q 686.97,217.32 690.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,210.00 Q 682.68,206.97 676.80,210.00 Q 682.68,213.03 690.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,210.00 Q 686.97,202.68 680.67,200.67 Q 682.68,206.97 690.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,210.00 Q 693.03,202.68 690.00,196.80 Q 686.97,202.68 690.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,210.00 Q 697.32,206.97 699.33,200.67 Q 693.03,202.68 690.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,210.00 Q 690.93,213.48 695.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,210.00 Q 686.52,210.93 684.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,210.00 Q 689.07,206.52 684.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,210.00 Q 693.48,209.07 695.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="690.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 690.00,225.12 C 683.60,218.72 676.74,211.86 674.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,194.88 C 696.40,201.28 703.26,208.14 705.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 775.20,210.00 C 764.22,220.98 753.42,231.78 750.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 724.80,210.00 C 735.78,199.02 746.58,188.22 750.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,225.12 C 743.60,218.72 736.74,211.86 734.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,194.88 C 756.40,201.28 763.26,208.14 765.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 810.00,184.80 C 820.98,195.78 831.78,206.58 835.20,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,235.20 C 799.02,224.22 788.22,213.42 784.80,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 810.00,210.00 Q 817.32,213.03 823.20,210.00 Q 817.32,206.97 810.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,210.00 Q 813.03,217.32 819.33,219.33 Q 817.32,213.03 810.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,210.00 Q 806.97,217.32 810.00,223.20 Q 813.03,217.32 810.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,210.00 Q 802.68,213.03 800.67,219.33 Q 806.97,217.32 810.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,210.00 Q 802.68,206.97 796.80,210.00 Q 802.68,213.03 810.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,210.00 Q 806.97,202.68 800.67,200.67 Q 802.68,206.97 810.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,210.00 Q 813.03,202.68 810.00,196.80 Q 806.97,202.68 810.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,210.00 Q 817.32,206.97 819.33,200.67 Q 813.03,202.68 810.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,210.00 Q 810.93,213.48 815.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,210.00 Q 806.52,210.93 804.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,210.00 Q 809.07,206.52 804.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,210.00 Q 813.48,209.07 815.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="810.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 825.12,210.00 C 818.72,216.40 811.86,223.26 810.00,225.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 794.88,210.00 C 801.28,203.60 808.14,196.74 810.00,194.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 844.80,210.00 C 855.78,199.02 866.58,188.22 870.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 895.20,210.00 C 884.22,220.98 873.42,231.78 870.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,210.00 Q 877.32,213.03 883.20,210.00 Q 877.32,206.97 870.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,210.00 Q 873.03,217.32 879.33,219.33 Q 877.32,213.03 870.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,210.00 Q 866.97,217.32 870.00,223.20 Q 873.03,217.32 870.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,210.00 Q 862.68,213.03 860.67,219.33 Q 866.97,217.32 870.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,210.00 Q 862.68,206.97 856.80,210.00 Q 862.68,213.03 870.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,210.00 Q 866.97,202.68 860.67,200.67 Q 862.68,206.97 870.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,210.00 Q 873.03,202.68 870.00,196.80 Q 866.97,202.68 870.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,210.00 Q 877.32,206.97 879.33,200.67 Q 873.03,202.68 870.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,210.00 Q 870.93,213.48 875.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,210.00 Q 866.52,210.93 864.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,210.00 Q 869.07,206.52 864.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,210.00 Q 873.48,209.07 875.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 870.00,194.88 C 876.40,201.28 883.26,208.14 885.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,225.12 C 863.60,218.72 856.74,211.86 854.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 930.00,184.80 C 940.98,195.78 951.78,206.58 955.20,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,235.20 C 919.02,224.22 908.22,213.42 904.80,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 945.12,210.00 C 938.72,216.40 931.86,223.26 930.00,225.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 914.88,210.00 C 921.28,203.60 928.14,196.74 930.00,194.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,184.80 C 1000.98,195.78 1011.78,206.58 1015.20,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,235.20 C 979.02,224.22 968.22,213.42 964.80,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1005.12,210.00 C 998.72,216.40 991.86,223.26 990.00,225.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 974.88,210.00 C 981.28,203.60 988.14,196.74 990.00,194.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,210.00 C 1035.78,199.02 1046.58,188.22 1050.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,210.00 C 1064.22,220.98 1053.42,231.78 1050.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,194.88 C 1056.40,201.28 1063.26,208.14 1065.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,225.12 C 1043.60,218.72 1036.74,211.86 1034.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1084.80,210.00 C 1095.78,199.02 1106.58,188.22 1110.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1135.20,210.00 C 1124.22,220.98 1113.42,231.78 1110.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1110.00,210.00 Q 1117.32,213.03 1123.20,210.00 Q 1117.32,206.97 1110.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,210.00 Q 1113.03,217.32 1119.33,219.33 Q 1117.32,213.03 1110.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,210.00 Q 1106.97,217.32 1110.00,223.20 Q 1113.03,217.32 1110.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,210.00 Q 1102.68,213.03 1100.67,219.33 Q 1106.97,217.32 1110.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,210.00 Q 1102.68,206.97 1096.80,210.00 Q 1102.68,213.03 1110.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,210.00 Q 1106.97,202.68 1100.67,200.67 Q 1102.68,206.97 1110.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,210.00 Q 1113.03,202.68 1110.00,196.80 Q 1106.97,202.68 1110.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,210.00 Q 1117.32,206.97 1119.33,200.67 Q 1113.03,202.68 1110.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,210.00 Q 1110.93,213.48 1115.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,210.00 Q 1106.52,210.93 1104.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,210.00 Q 1109.07,206.52 1104.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,210.00 Q 1113.48,209.07 1115.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1110.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1110.00,194.88 C 1116.40,201.28 1123.26,208.14 1125.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,225.12 C 1103.60,218.72 1096.74,211.86 1094.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1195.20,210.00 C 1184.22,220.98 1173.42,231.78 1170.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1144.80,210.00 C 1155.78,199.02 1166.58,188.22 1170.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1170.00,225.12 C 1163.60,218.72 1156.74,211.86 1154.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,194.88 C 1176.40,201.28 1183.26,208.14 1185.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1255.20,210.00 C 1244.22,220.98 1233.42,231.78 1230.00,235.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1204.80,210.00 C 1215.78,199.02 1226.58,188.22 1230.00,184.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1230.00,225.12 C 1223.60,218.72 1216.74,211.86 1214.88,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,194.88 C 1236.40,201.28 1243.26,208.14 1245.12,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1290.00,184.80 C 1300.98,195.78 1311.78,206.58 1315.20,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,235.20 C 1279.02,224.22 1268.22,213.42 1264.80,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1290.00,210.00 Q 1297.32,213.03 1303.20,210.00 Q 1297.32,206.97 1290.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,210.00 Q 1293.03,217.32 1299.33,219.33 Q 1297.32,213.03 1290.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,210.00 Q 1286.97,217.32 1290.00,223.20 Q 1293.03,217.32 1290.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,210.00 Q 1282.68,213.03 1280.67,219.33 Q 1286.97,217.32 1290.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,210.00 Q 1282.68,206.97 1276.80,210.00 Q 1282.68,213.03 1290.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,210.00 Q 1286.97,202.68 1280.67,200.67 Q 1282.68,206.97 1290.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,210.00 Q 1293.03,202.68 1290.00,196.80 Q 1286.97,202.68 1290.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,210.00 Q 1297.32,206.97 1299.33,200.67 Q 1293.03,202.68 1290.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,210.00 Q 1290.93,213.48 1295.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,210.00 Q 1286.52,210.93 1284.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,210.00 Q 1289.07,206.52 1284.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,210.00 Q 1293.48,209.07 1295.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1290.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1305.12,210.00 C 1298.72,216.40 1291.86,223.26 1290.00,225.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1274.88,210.00 C 1281.28,203.60 1288.14,196.74 1290.00,194.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1350.00,184.80 C 1360.98,195.78 1371.78,206.58 1375.20,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,235.20 C 1339.02,224.22 1328.22,213.42 1324.80,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1350.00,210.00 Q 1357.32,213.03 1363.20,210.00 Q 1357.32,206.97 1350.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,210.00 Q 1353.03,217.32 1359.33,219.33 Q 1357.32,213.03 1350.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,210.00 Q 1346.97,217.32 1350.00,223.20 Q 1353.03,217.32 1350.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,210.00 Q 1342.68,213.03 1340.67,219.33 Q 1346.97,217.32 1350.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,210.00 Q 1342.68,206.97 1336.80,210.00 Q 1342.68,213.03 1350.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,210.00 Q 1346.97,202.68 1340.67,200.67 Q 1342.68,206.97 1350.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,210.00 Q 1353.03,202.68 1350.00,196.80 Q 1346.97,202.68 1350.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,210.00 Q 1357.32,206.97 1359.33,200.67 Q 1353.03,202.68 1350.00,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,210.00 Q 1350.93,213.48 1355.09,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,210.00 Q 1346.52,210.93 1344.91,215.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,210.00 Q 1349.07,206.52 1344.91,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,210.00 Q 1353.48,209.07 1355.09,204.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1350.0" cy="210.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1365.12,210.00 C 1358.72,216.40 1351.86,223.26 1350.00,225.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1334.88,210.00 C 1341.28,203.60 1348.14,196.74 1350.00,194.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,295.20 C 139.02,284.22 128.22,273.42 124.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,244.80 C 160.98,255.78 171.78,266.58 175.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 134.88,270.00 C 141.28,263.60 148.14,256.74 150.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 165.12,270.00 C 158.72,276.40 151.86,283.26 150.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 210.00,295.20 C 199.02,284.22 188.22,273.42 184.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,244.80 C 220.98,255.78 231.78,266.58 235.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 210.00,270.00 Q 217.32,273.03 223.20,270.00 Q 217.32,266.97 210.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,270.00 Q 213.03,277.32 219.33,279.33 Q 217.32,273.03 210.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,270.00 Q 206.97,277.32 210.00,283.20 Q 213.03,277.32 210.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,270.00 Q 202.68,273.03 200.67,279.33 Q 206.97,277.32 210.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,270.00 Q 202.68,266.97 196.80,270.00 Q 202.68,273.03 210.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,270.00 Q 206.97,262.68 200.67,260.67 Q 202.68,266.97 210.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,270.00 Q 213.03,262.68 210.00,256.80 Q 206.97,262.68 210.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,270.00 Q 217.32,266.97 219.33,260.67 Q 213.03,262.68 210.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,270.00 Q 210.93,273.48 215.09,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,270.00 Q 206.52,270.93 204.91,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,270.00 Q 209.07,266.52 204.91,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,270.00 Q 213.48,269.07 215.09,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="210.0" cy="270.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 194.88,270.00 C 201.28,263.60 208.14,256.74 210.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 225.12,270.00 C 218.72,276.40 211.86,283.26 210.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,244.80 C 280.98,255.78 291.78,266.58 295.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,295.20 C 259.02,284.22 248.22,273.42 244.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 285.12,270.00 C 278.72,276.40 271.86,283.26 270.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 254.88,270.00 C 261.28,263.60 268.14,256.74 270.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,270.00 C 315.78,259.02 326.58,248.22 330.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,270.00 C 344.22,280.98 333.42,291.78 330.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 330.00,270.00 Q 337.32,273.03 343.20,270.00 Q 337.32,266.97 330.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,270.00 Q 333.03,277.32 339.33,279.33 Q 337.32,273.03 330.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,270.00 Q 326.97,277.32 330.00,283.20 Q 333.03,277.32 330.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,270.00 Q 322.68,273.03 320.67,279.33 Q 326.97,277.32 330.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,270.00 Q 322.68,266.97 316.80,270.00 Q 322.68,273.03 330.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,270.00 Q 326.97,262.68 320.67,260.67 Q 322.68,266.97 330.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,270.00 Q 333.03,262.68 330.00,256.80 Q 326.97,262.68 330.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,270.00 Q 337.32,266.97 339.33,260.67 Q 333.03,262.68 330.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,270.00 Q 330.93,273.48 335.09,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,270.00 Q 326.52,270.93 324.91,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,270.00 Q 329.07,266.52 324.91,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,270.00 Q 333.48,269.07 335.09,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="330.0" cy="270.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 330.00,254.88 C 336.40,261.28 343.26,268.14 345.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,285.12 C 323.60,278.72 316.74,271.86 314.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 390.00,295.20 C 379.02,284.22 368.22,273.42 364.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,244.80 C 400.98,255.78 411.78,266.58 415.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 374.88,270.00 C 381.28,263.60 388.14,256.74 390.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 405.12,270.00 C 398.72,276.40 391.86,283.26 390.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 450.00,244.80 C 460.98,255.78 471.78,266.58 475.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,295.20 C 439.02,284.22 428.22,273.42 424.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 450.00,270.00 Q 457.32,273.03 463.20,270.00 Q 457.32,266.97 450.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,270.00 Q 453.03,277.32 459.33,279.33 Q 457.32,273.03 450.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,270.00 Q 446.97,277.32 450.00,283.20 Q 453.03,277.32 450.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,270.00 Q 442.68,273.03 440.67,279.33 Q 446.97,277.32 450.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,270.00 Q 442.68,266.97 436.80,270.00 Q 442.68,273.03 450.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,270.00 Q 446.97,262.68 440.67,260.67 Q 442.68,266.97 450.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,270.00 Q 453.03,262.68 450.00,256.80 Q 446.97,262.68 450.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,270.00 Q 457.32,266.97 459.33,260.67 Q 453.03,262.68 450.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,270.00 Q 450.93,273.48 455.09,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,270.00 Q 446.52,270.93 444.91,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,270.00 Q 449.07,266.52 444.91,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,270.00 Q 453.48,269.07 455.09,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="450.0" cy="270.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 465.12,270.00 C 458.72,276.40 451.86,283.26 450.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 434.88,270.00 C 441.28,263.60 448.14,256.74 450.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 484.80,270.00 C 495.78,259.02 506.58,248.22 510.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 535.20,270.00 C 524.22,280.98 513.42,291.78 510.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,270.00 Q 517.32,273.03 523.20,270.00 Q 517.32,266.97 510.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,270.00 Q 513.03,277.32 519.33,279.33 Q 517.32,273.03 510.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,270.00 Q 506.97,277.32 510.00,283.20 Q 513.03,277.32 510.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,270.00 Q 502.68,273.03 500.67,279.33 Q 506.97,277.32 510.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,270.00 Q 502.68,266.97 496.80,270.00 Q 502.68,273.03 510.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,270.00 Q 506.97,262.68 500.67,260.67 Q 502.68,266.97 510.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,270.00 Q 513.03,262.68 510.00,256.80 Q 506.97,262.68 510.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,270.00 Q 517.32,266.97 519.33,260.67 Q 513.03,262.68 510.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,270.00 Q 510.93,273.48 515.09,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,270.00 Q 506.52,270.93 504.91,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,270.00 Q 509.07,266.52 504.91,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,270.00 Q 513.48,269.07 515.09,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="270.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 510.00,254.88 C 516.40,261.28 523.26,268.14 525.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,285.12 C 503.60,278.72 496.74,271.86 494.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,270.00 C 555.78,259.02 566.58,248.22 570.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,270.00 C 584.22,280.98 573.42,291.78 570.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 570.00,254.88 C 576.40,261.28 583.26,268.14 585.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,285.12 C 563.60,278.72 556.74,271.86 554.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,270.00 C 615.78,259.02 626.58,248.22 630.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,270.00 C 644.22,280.98 633.42,291.78 630.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,254.88 C 636.40,261.28 643.26,268.14 645.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,285.12 C 623.60,278.72 616.74,271.86 614.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 690.00,295.20 C 679.02,284.22 668.22,273.42 664.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,244.80 C 700.98,255.78 711.78,266.58 715.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 690.00,270.00 Q 697.32,273.03 703.20,270.00 Q 697.32,266.97 690.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,270.00 Q 693.03,277.32 699.33,279.33 Q 697.32,273.03 690.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,270.00 Q 686.97,277.32 690.00,283.20 Q 693.03,277.32 690.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,270.00 Q 682.68,273.03 680.67,279.33 Q 686.97,277.32 690.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,270.00 Q 682.68,266.97 676.80,270.00 Q 682.68,273.03 690.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,270.00 Q 686.97,262.68 680.67,260.67 Q 682.68,266.97 690.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,270.00 Q 693.03,262.68 690.00,256.80 Q 686.97,262.68 690.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,270.00 Q 697.32,266.97 699.33,260.67 Q 693.03,262.68 690.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,270.00 Q 690.93,273.48 695.09,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,270.00 Q 686.52,270.93 684.91,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,270.00 Q 689.07,266.52 684.91,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,270.00 Q 693.48,269.07 695.09,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="690.0" cy="270.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 674.88,270.00 C 681.28,263.60 688.14,256.74 690.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 705.12,270.00 C 698.72,276.40 691.86,283.26 690.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 750.00,244.80 C 760.98,255.78 771.78,266.58 775.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,295.20 C 739.02,284.22 728.22,273.42 724.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 765.12,270.00 C 758.72,276.40 751.86,283.26 750.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 734.88,270.00 C 741.28,263.60 748.14,256.74 750.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 784.80,270.00 C 795.78,259.02 806.58,248.22 810.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 835.20,270.00 C 824.22,280.98 813.42,291.78 810.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 810.00,270.00 Q 817.32,273.03 823.20,270.00 Q 817.32,266.97 810.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,270.00 Q 813.03,277.32 819.33,279.33 Q 817.32,273.03 810.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,270.00 Q 806.97,277.32 810.00,283.20 Q 813.03,277.32 810.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,270.00 Q 802.68,273.03 800.67,279.33 Q 806.97,277.32 810.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,270.00 Q 802.68,266.97 796.80,270.00 Q 802.68,273.03 810.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,270.00 Q 806.97,262.68 800.67,260.67 Q 802.68,266.97 810.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,270.00 Q 813.03,262.68 810.00,256.80 Q 806.97,262.68 810.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,270.00 Q 817.32,266.97 819.33,260.67 Q 813.03,262.68 810.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,270.00 Q 810.93,273.48 815.09,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,270.00 Q 806.52,270.93 804.91,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,270.00 Q 809.07,266.52 804.91,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,270.00 Q 813.48,269.07 815.09,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="810.0" cy="270.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 810.00,254.88 C 816.40,261.28 823.26,268.14 825.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,285.12 C 803.60,278.72 796.74,271.86 794.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 895.20,270.00 C 884.22,280.98 873.42,291.78 870.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 844.80,270.00 C 855.78,259.02 866.58,248.22 870.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 870.00,285.12 C 863.60,278.72 856.74,271.86 854.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,254.88 C 876.40,261.28 883.26,268.14 885.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 955.20,270.00 C 944.22,280.98 933.42,291.78 930.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 904.80,270.00 C 915.78,259.02 926.58,248.22 930.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,270.00 Q 937.32,273.03 943.20,270.00 Q 937.32,266.97 930.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,270.00 Q 933.03,277.32 939.33,279.33 Q 937.32,273.03 930.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,270.00 Q 926.97,277.32 930.00,283.20 Q 933.03,277.32 930.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,270.00 Q 922.68,273.03 920.67,279.33 Q 926.97,277.32 930.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,270.00 Q 922.68,266.97 916.80,270.00 Q 922.68,273.03 930.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,270.00 Q 926.97,262.68 920.67,260.67 Q 922.68,266.97 930.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,270.00 Q 933.03,262.68 930.00,256.80 Q 926.97,262.68 930.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,270.00 Q 937.32,266.97 939.33,260.67 Q 933.03,262.68 930.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,270.00 Q 930.93,273.48 935.09,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,270.00 Q 926.52,270.93 924.91,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,270.00 Q 929.07,266.52 924.91,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,270.00 Q 933.48,269.07 935.09,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="270.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 930.00,285.12 C 923.60,278.72 916.74,271.86 914.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,254.88 C 936.40,261.28 943.26,268.14 945.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,244.80 C 1000.98,255.78 1011.78,266.58 1015.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,295.20 C 979.02,284.22 968.22,273.42 964.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 990.00,270.00 Q 997.32,273.03 1003.20,270.00 Q 997.32,266.97 990.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,270.00 Q 993.03,277.32 999.33,279.33 Q 997.32,273.03 990.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,270.00 Q 986.97,277.32 990.00,283.20 Q 993.03,277.32 990.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,270.00 Q 982.68,273.03 980.67,279.33 Q 986.97,277.32 990.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,270.00 Q 982.68,266.97 976.80,270.00 Q 982.68,273.03 990.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,270.00 Q 986.97,262.68 980.67,260.67 Q 982.68,266.97 990.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,270.00 Q 993.03,262.68 990.00,256.80 Q 986.97,262.68 990.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,270.00 Q 997.32,266.97 999.33,260.67 Q 993.03,262.68 990.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,270.00 Q 990.93,273.48 995.09,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,270.00 Q 986.52,270.93 984.91,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,270.00 Q 989.07,266.52 984.91,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,270.00 Q 993.48,269.07 995.09,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="990.0" cy="270.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1005.12,270.00 C 998.72,276.40 991.86,283.26 990.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 974.88,270.00 C 981.28,263.60 988.14,256.74 990.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1075.20,270.00 C 1064.22,280.98 1053.42,291.78 1050.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1024.80,270.00 C 1035.78,259.02 1046.58,248.22 1050.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,285.12 C 1043.60,278.72 1036.74,271.86 1034.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,254.88 C 1056.40,261.28 1063.26,268.14 1065.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1110.00,295.20 C 1099.02,284.22 1088.22,273.42 1084.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,244.80 C 1120.98,255.78 1131.78,266.58 1135.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1094.88,270.00 C 1101.28,263.60 1108.14,256.74 1110.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1125.12,270.00 C 1118.72,276.40 1111.86,283.26 1110.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1170.00,295.20 C 1159.02,284.22 1148.22,273.42 1144.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,244.80 C 1180.98,255.78 1191.78,266.58 1195.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1170.00,270.00 Q 1177.32,273.03 1183.20,270.00 Q 1177.32,266.97 1170.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,270.00 Q 1173.03,277.32 1179.33,279.33 Q 1177.32,273.03 1170.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,270.00 Q 1166.97,277.32 1170.00,283.20 Q 1173.03,277.32 1170.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,270.00 Q 1162.68,273.03 1160.67,279.33 Q 1166.97,277.32 1170.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,270.00 Q 1162.68,266.97 1156.80,270.00 Q 1162.68,273.03 1170.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,270.00 Q 1166.97,262.68 1160.67,260.67 Q 1162.68,266.97 1170.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,270.00 Q 1173.03,262.68 1170.00,256.80 Q 1166.97,262.68 1170.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,270.00 Q 1177.32,266.97 1179.33,260.67 Q 1173.03,262.68 1170.00,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,270.00 Q 1170.93,273.48 1175.09,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,270.00 Q 1166.52,270.93 1164.91,275.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,270.00 Q 1169.07,266.52 1164.91,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,270.00 Q 1173.48,269.07 1175.09,264.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1170.0" cy="270.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1154.88,270.00 C 1161.28,263.60 1168.14,256.74 1170.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1185.12,270.00 C 1178.72,276.40 1171.86,283.26 1170.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,244.80 C 1240.98,255.78 1251.78,266.58 1255.20,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,295.20 C 1219.02,284.22 1208.22,273.42 1204.80,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1245.12,270.00 C 1238.72,276.40 1231.86,283.26 1230.00,285.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1214.88,270.00 C 1221.28,263.60 1228.14,256.74 1230.00,254.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1264.80,270.00 C 1275.78,259.02 1286.58,248.22 1290.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1315.20,270.00 C 1304.22,280.98 1293.42,291.78 1290.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1290.00,254.88 C 1296.40,261.28 1303.26,268.14 1305.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,285.12 C 1283.60,278.72 1276.74,271.86 1274.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1375.20,270.00 C 1364.22,280.98 1353.42,291.78 1350.00,295.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1324.80,270.00 C 1335.78,259.02 1346.58,248.22 1350.00,244.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,285.12 C 1343.60,278.72 1336.74,271.86 1334.88,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,254.88 C 1356.40,261.28 1363.26,268.14 1365.12,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 124.80,330.00 C 135.78,319.02 146.58,308.22 150.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 175.20,330.00 C 164.22,340.98 153.42,351.78 150.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 150.00,314.88 C 156.40,321.28 163.26,328.14 165.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,345.12 C 143.60,338.72 136.74,331.86 134.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 210.00,304.80 C 220.98,315.78 231.78,326.58 235.20,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,355.20 C 199.02,344.22 188.22,333.42 184.80,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 210.00,330.00 Q 217.32,333.03 223.20,330.00 Q 217.32,326.97 210.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,330.00 Q 213.03,337.32 219.33,339.33 Q 217.32,333.03 210.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,330.00 Q 206.97,337.32 210.00,343.20 Q 213.03,337.32 210.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,330.00 Q 202.68,333.03 200.67,339.33 Q 206.97,337.32 210.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,330.00 Q 202.68,326.97 196.80,330.00 Q 202.68,333.03 210.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,330.00 Q 206.97,322.68 200.67,320.67 Q 202.68,326.97 210.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,330.00 Q 213.03,322.68 210.00,316.80 Q 206.97,322.68 210.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,330.00 Q 217.32,326.97 219.33,320.67 Q 213.03,322.68 210.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,330.00 Q 210.93,333.48 215.09,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,330.00 Q 206.52,330.93 204.91,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,330.00 Q 209.07,326.52 204.91,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,330.00 Q 213.48,329.07 215.09,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="210.0" cy="330.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 225.12,330.00 C 218.72,336.40 211.86,343.26 210.00,345.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 194.88,330.00 C 201.28,323.60 208.14,316.74 210.00,314.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 295.20,330.00 C 284.22,340.98 273.42,351.78 270.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 244.80,330.00 C 255.78,319.02 266.58,308.22 270.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 270.00,345.12 C 263.60,338.72 256.74,331.86 254.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,314.88 C 276.40,321.28 283.26,328.14 285.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 330.00,355.20 C 319.02,344.22 308.22,333.42 304.80,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,304.80 C 340.98,315.78 351.78,326.58 355.20,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 314.88,330.00 C 321.28,323.60 328.14,316.74 330.00,314.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 345.12,330.00 C 338.72,336.40 331.86,343.26 330.00,345.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 390.00,355.20 C 379.02,344.22 368.22,333.42 364.80,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,304.80 C 400.98,315.78 411.78,326.58 415.20,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 374.88,330.00 C 381.28,323.60 388.14,316.74 390.00,314.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 405.12,330.00 C 398.72,336.40 391.86,343.26 390.00,345.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 475.20,330.00 C 464.22,340.98 453.42,351.78 450.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 424.80,330.00 C 435.78,319.02 446.58,308.22 450.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 450.00,330.00 Q 457.32,333.03 463.20,330.00 Q 457.32,326.97 450.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,330.00 Q 453.03,337.32 459.33,339.33 Q 457.32,333.03 450.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,330.00 Q 446.97,337.32 450.00,343.20 Q 453.03,337.32 450.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,330.00 Q 442.68,333.03 440.67,339.33 Q 446.97,337.32 450.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,330.00 Q 442.68,326.97 436.80,330.00 Q 442.68,333.03 450.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,330.00 Q 446.97,322.68 440.67,320.67 Q 442.68,326.97 450.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,330.00 Q 453.03,322.68 450.00,316.80 Q 446.97,322.68 450.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,330.00 Q 457.32,326.97 459.33,320.67 Q 453.03,322.68 450.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,330.00 Q 450.93,333.48 455.09,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,330.00 Q 446.52,330.93 444.91,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,330.00 Q 449.07,326.52 444.91,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,330.00 Q 453.48,329.07 455.09,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="450.0" cy="330.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 450.00,345.12 C 443.60,338.72 436.74,331.86 434.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,314.88 C 456.40,321.28 463.26,328.14 465.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 484.80,330.00 C 495.78,319.02 506.58,308.22 510.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 535.20,330.00 C 524.22,340.98 513.42,351.78 510.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,330.00 Q 517.32,333.03 523.20,330.00 Q 517.32,326.97 510.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,330.00 Q 513.03,337.32 519.33,339.33 Q 517.32,333.03 510.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,330.00 Q 506.97,337.32 510.00,343.20 Q 513.03,337.32 510.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,330.00 Q 502.68,333.03 500.67,339.33 Q 506.97,337.32 510.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,330.00 Q 502.68,326.97 496.80,330.00 Q 502.68,333.03 510.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,330.00 Q 506.97,322.68 500.67,320.67 Q 502.68,326.97 510.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,330.00 Q 513.03,322.68 510.00,316.80 Q 506.97,322.68 510.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,330.00 Q 517.32,326.97 519.33,320.67 Q 513.03,322.68 510.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,330.00 Q 510.93,333.48 515.09,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,330.00 Q 506.52,330.93 504.91,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,330.00 Q 509.07,326.52 504.91,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,330.00 Q 513.48,329.07 515.09,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="330.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 510.00,314.88 C 516.40,321.28 523.26,328.14 525.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,345.12 C 503.60,338.72 496.74,331.86 494.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 595.20,330.00 C 584.22,340.98 573.42,351.78 570.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 544.80,330.00 C 555.78,319.02 566.58,308.22 570.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 570.00,345.12 C 563.60,338.72 556.74,331.86 554.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,314.88 C 576.40,321.28 583.26,328.14 585.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 655.20,330.00 C 644.22,340.98 633.42,351.78 630.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 604.80,330.00 C 615.78,319.02 626.58,308.22 630.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,345.12 C 623.60,338.72 616.74,331.86 614.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,314.88 C 636.40,321.28 643.26,328.14 645.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 690.00,304.80 C 700.98,315.78 711.78,326.58 715.20,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,355.20 C 679.02,344.22 668.22,333.42 664.80,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 690.00,330.00 Q 697.32,333.03 703.20,330.00 Q 697.32,326.97 690.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,330.00 Q 693.03,337.32 699.33,339.33 Q 697.32,333.03 690.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,330.00 Q 686.97,337.32 690.00,343.20 Q 693.03,337.32 690.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,330.00 Q 682.68,333.03 680.67,339.33 Q 686.97,337.32 690.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,330.00 Q 682.68,326.97 676.80,330.00 Q 682.68,333.03 690.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,330.00 Q 686.97,322.68 680.67,320.67 Q 682.68,326.97 690.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,330.00 Q 693.03,322.68 690.00,316.80 Q 686.97,322.68 690.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,330.00 Q 697.32,326.97 699.33,320.67 Q 693.03,322.68 690.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,330.00 Q 690.93,333.48 695.09,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,330.00 Q 686.52,330.93 684.91,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,330.00 Q 689.07,326.52 684.91,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,330.00 Q 693.48,329.07 695.09,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="690.0" cy="330.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 705.12,330.00 C 698.72,336.40 691.86,343.26 690.00,345.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 674.88,330.00 C 681.28,323.60 688.14,316.74 690.00,314.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 750.00,304.80 C 760.98,315.78 771.78,326.58 775.20,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,355.20 C 739.02,344.22 728.22,333.42 724.80,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 750.00,330.00 Q 757.32,333.03 763.20,330.00 Q 757.32,326.97 750.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,330.00 Q 753.03,337.32 759.33,339.33 Q 757.32,333.03 750.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,330.00 Q 746.97,337.32 750.00,343.20 Q 753.03,337.32 750.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,330.00 Q 742.68,333.03 740.67,339.33 Q 746.97,337.32 750.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,330.00 Q 742.68,326.97 736.80,330.00 Q 742.68,333.03 750.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,330.00 Q 746.97,322.68 740.67,320.67 Q 742.68,326.97 750.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,330.00 Q 753.03,322.68 750.00,316.80 Q 746.97,322.68 750.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,330.00 Q 757.32,326.97 759.33,320.67 Q 753.03,322.68 750.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,330.00 Q 750.93,333.48 755.09,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,330.00 Q 746.52,330.93 744.91,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,330.00 Q 749.07,326.52 744.91,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,330.00 Q 753.48,329.07 755.09,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="750.0" cy="330.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 765.12,330.00 C 758.72,336.40 751.86,343.26 750.00,345.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 734.88,330.00 C 741.28,323.60 748.14,316.74 750.00,314.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 835.20,330.00 C 824.22,340.98 813.42,351.78 810.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 784.80,330.00 C 795.78,319.02 806.58,308.22 810.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,345.12 C 803.60,338.72 796.74,331.86 794.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,314.88 C 816.40,321.28 823.26,328.14 825.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 870.00,355.20 C 859.02,344.22 848.22,333.42 844.80,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,304.80 C 880.98,315.78 891.78,326.58 895.20,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 854.88,330.00 C 861.28,323.60 868.14,316.74 870.00,314.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 885.12,330.00 C 878.72,336.40 871.86,343.26 870.00,345.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 904.80,330.00 C 915.78,319.02 926.58,308.22 930.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 955.20,330.00 C 944.22,340.98 933.42,351.78 930.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,330.00 Q 937.32,333.03 943.20,330.00 Q 937.32,326.97 930.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,330.00 Q 933.03,337.32 939.33,339.33 Q 937.32,333.03 930.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,330.00 Q 926.97,337.32 930.00,343.20 Q 933.03,337.32 930.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,330.00 Q 922.68,333.03 920.67,339.33 Q 926.97,337.32 930.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,330.00 Q 922.68,326.97 916.80,330.00 Q 922.68,333.03 930.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,330.00 Q 926.97,322.68 920.67,320.67 Q 922.68,326.97 930.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,330.00 Q 933.03,322.68 930.00,316.80 Q 926.97,322.68 930.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,330.00 Q 937.32,326.97 939.33,320.67 Q 933.03,322.68 930.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,330.00 Q 930.93,333.48 935.09,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,330.00 Q 926.52,330.93 924.91,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,330.00 Q 929.07,326.52 924.91,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,330.00 Q 933.48,329.07 935.09,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="330.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 930.00,314.88 C 936.40,321.28 943.26,328.14 945.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,345.12 C 923.60,338.72 916.74,331.86 914.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1015.20,330.00 C 1004.22,340.98 993.42,351.78 990.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 964.80,330.00 C 975.78,319.02 986.58,308.22 990.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 990.00,345.12 C 983.60,338.72 976.74,331.86 974.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,314.88 C 996.40,321.28 1003.26,328.14 1005.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1075.20,330.00 C 1064.22,340.98 1053.42,351.78 1050.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1024.80,330.00 C 1035.78,319.02 1046.58,308.22 1050.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,345.12 C 1043.60,338.72 1036.74,331.86 1034.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,314.88 C 1056.40,321.28 1063.26,328.14 1065.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1084.80,330.00 C 1095.78,319.02 1106.58,308.22 1110.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1135.20,330.00 C 1124.22,340.98 1113.42,351.78 1110.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1110.00,314.88 C 1116.40,321.28 1123.26,328.14 1125.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,345.12 C 1103.60,338.72 1096.74,331.86 1094.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1170.00,304.80 C 1180.98,315.78 1191.78,326.58 1195.20,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,355.20 C 1159.02,344.22 1148.22,333.42 1144.80,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1170.00,330.00 Q 1177.32,333.03 1183.20,330.00 Q 1177.32,326.97 1170.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,330.00 Q 1173.03,337.32 1179.33,339.33 Q 1177.32,333.03 1170.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,330.00 Q 1166.97,337.32 1170.00,343.20 Q 1173.03,337.32 1170.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,330.00 Q 1162.68,333.03 1160.67,339.33 Q 1166.97,337.32 1170.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,330.00 Q 1162.68,326.97 1156.80,330.00 Q 1162.68,333.03 1170.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,330.00 Q 1166.97,322.68 1160.67,320.67 Q 1162.68,326.97 1170.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,330.00 Q 1173.03,322.68 1170.00,316.80 Q 1166.97,322.68 1170.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,330.00 Q 1177.32,326.97 1179.33,320.67 Q 1173.03,322.68 1170.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,330.00 Q 1170.93,333.48 1175.09,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,330.00 Q 1166.52,330.93 1164.91,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,330.00 Q 1169.07,326.52 1164.91,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,330.00 Q 1173.48,329.07 1175.09,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1170.0" cy="330.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1185.12,330.00 C 1178.72,336.40 1171.86,343.26 1170.00,345.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1154.88,330.00 C 1161.28,323.60 1168.14,316.74 1170.00,314.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1204.80,330.00 C 1215.78,319.02 1226.58,308.22 1230.00,304.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1255.20,330.00 C 1244.22,340.98 1233.42,351.78 1230.00,355.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1230.00,330.00 Q 1237.32,333.03 1243.20,330.00 Q 1237.32,326.97 1230.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,330.00 Q 1233.03,337.32 1239.33,339.33 Q 1237.32,333.03 1230.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,330.00 Q 1226.97,337.32 1230.00,343.20 Q 1233.03,337.32 1230.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,330.00 Q 1222.68,333.03 1220.67,339.33 Q 1226.97,337.32 1230.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,330.00 Q 1222.68,326.97 1216.80,330.00 Q 1222.68,333.03 1230.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,330.00 Q 1226.97,322.68 1220.67,320.67 Q 1222.68,326.97 1230.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,330.00 Q 1233.03,322.68 1230.00,316.80 Q 1226.97,322.68 1230.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,330.00 Q 1237.32,326.97 1239.33,320.67 Q 1233.03,322.68 1230.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,330.00 Q 1230.93,333.48 1235.09,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,330.00 Q 1226.52,330.93 1224.91,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,330.00 Q 1229.07,326.52 1224.91,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,330.00 Q 1233.48,329.07 1235.09,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1230.0" cy="330.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1230.00,314.88 C 1236.40,321.28 1243.26,328.14 1245.12,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,345.12 C 1223.60,338.72 1216.74,331.86 1214.88,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1290.00,304.80 C 1300.98,315.78 1311.78,326.58 1315.20,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,355.20 C 1279.02,344.22 1268.22,333.42 1264.80,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1305.12,330.00 C 1298.72,336.40 1291.86,343.26 1290.00,345.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1274.88,330.00 C 1281.28,323.60 1288.14,316.74 1290.00,314.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1350.00,355.20 C 1339.02,344.22 1328.22,333.42 1324.80,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,304.80 C 1360.98,315.78 1371.78,326.58 1375.20,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1350.00,330.00 Q 1357.32,333.03 1363.20,330.00 Q 1357.32,326.97 1350.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,330.00 Q 1353.03,337.32 1359.33,339.33 Q 1357.32,333.03 1350.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,330.00 Q 1346.97,337.32 1350.00,343.20 Q 1353.03,337.32 1350.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,330.00 Q 1342.68,333.03 1340.67,339.33 Q 1346.97,337.32 1350.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,330.00 Q 1342.68,326.97 1336.80,330.00 Q 1342.68,333.03 1350.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,330.00 Q 1346.97,322.68 1340.67,320.67 Q 1342.68,326.97 1350.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,330.00 Q 1353.03,322.68 1350.00,316.80 Q 1346.97,322.68 1350.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,330.00 Q 1357.32,326.97 1359.33,320.67 Q 1353.03,322.68 1350.00,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,330.00 Q 1350.93,333.48 1355.09,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,330.00 Q 1346.52,330.93 1344.91,335.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,330.00 Q 1349.07,326.52 1344.91,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,330.00 Q 1353.48,329.07 1355.09,324.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1350.0" cy="330.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1334.88,330.00 C 1341.28,323.60 1348.14,316.74 1350.00,314.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1365.12,330.00 C 1358.72,336.40 1351.86,343.26 1350.00,345.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,364.80 C 160.98,375.78 171.78,386.58 175.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,415.20 C 139.02,404.22 128.22,393.42 124.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,390.00 Q 157.32,393.03 163.20,390.00 Q 157.32,386.97 150.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,390.00 Q 153.03,397.32 159.33,399.33 Q 157.32,393.03 150.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,390.00 Q 146.97,397.32 150.00,403.20 Q 153.03,397.32 150.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,390.00 Q 142.68,393.03 140.67,399.33 Q 146.97,397.32 150.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,390.00 Q 142.68,386.97 136.80,390.00 Q 142.68,393.03 150.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,390.00 Q 146.97,382.68 140.67,380.67 Q 142.68,386.97 150.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,390.00 Q 153.03,382.68 150.00,376.80 Q 146.97,382.68 150.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,390.00 Q 157.32,386.97 159.33,380.67 Q 153.03,382.68 150.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,390.00 Q 150.93,393.48 155.09,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,390.00 Q 146.52,390.93 144.91,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,390.00 Q 149.07,386.52 144.91,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,390.00 Q 153.48,389.07 155.09,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="390.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 165.12,390.00 C 158.72,396.40 151.86,403.26 150.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 134.88,390.00 C 141.28,383.60 148.14,376.74 150.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 235.20,390.00 C 224.22,400.98 213.42,411.78 210.00,415.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 184.80,390.00 C 195.78,379.02 206.58,368.22 210.00,364.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,405.12 C 203.60,398.72 196.74,391.86 194.88,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,374.88 C 216.40,381.28 223.26,388.14 225.12,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 295.20,390.00 C 284.22,400.98 273.42,411.78 270.00,415.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 244.80,390.00 C 255.78,379.02 266.58,368.22 270.00,364.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 270.00,405.12 C 263.60,398.72 256.74,391.86 254.88,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,374.88 C 276.40,381.28 283.26,388.14 285.12,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,390.00 C 315.78,379.02 326.58,368.22 330.00,364.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,390.00 C 344.22,400.98 333.42,411.78 330.00,415.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 330.00,374.88 C 336.40,381.28 343.26,388.14 345.12,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,405.12 C 323.60,398.72 316.74,391.86 314.88,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 390.00,364.80 C 400.98,375.78 411.78,386.58 415.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,415.20 C 379.02,404.22 368.22,393.42 364.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 390.00,390.00 Q 397.32,393.03 403.20,390.00 Q 397.32,386.97 390.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,390.00 Q 393.03,397.32 399.33,399.33 Q 397.32,393.03 390.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,390.00 Q 386.97,397.32 390.00,403.20 Q 393.03,397.32 390.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,390.00 Q 382.68,393.03 380.67,399.33 Q 386.97,397.32 390.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,390.00 Q 382.68,386.97 376.80,390.00 Q 382.68,393.03 390.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,390.00 Q 386.97,382.68 380.67,380.67 Q 382.68,386.97 390.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,390.00 Q 393.03,382.68 390.00,376.80 Q 386.97,382.68 390.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,390.00 Q 397.32,386.97 399.33,380.67 Q 393.03,382.68 390.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,390.00 Q 390.93,393.48 395.09,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,390.00 Q 386.52,390.93 384.91,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,390.00 Q 389.07,386.52 384.91,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,390.00 Q 393.48,389.07 395.09,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="390.0" cy="390.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 405.12,390.00 C 398.72,396.40 391.86,403.26 390.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 374.88,390.00 C 381.28,383.60 388.14,376.74 390.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 450.00,364.80 C 460.98,375.78 471.78,386.58 475.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,415.20 C 439.02,404.22 428.22,393.42 424.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 465.12,390.00 C 458.72,396.40 451.86,403.26 450.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 434.88,390.00 C 441.28,383.60 448.14,376.74 450.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,364.80 C 520.98,375.78 531.78,386.58 535.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,415.20 C 499.02,404.22 488.22,393.42 484.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 525.12,390.00 C 518.72,396.40 511.86,403.26 510.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 494.88,390.00 C 501.28,383.60 508.14,376.74 510.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 570.00,415.20 C 559.02,404.22 548.22,393.42 544.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,364.80 C 580.98,375.78 591.78,386.58 595.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 554.88,390.00 C 561.28,383.60 568.14,376.74 570.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 585.12,390.00 C 578.72,396.40 571.86,403.26 570.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 655.20,390.00 C 644.22,400.98 633.42,411.78 630.00,415.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 604.80,390.00 C 615.78,379.02 626.58,368.22 630.00,364.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 630.00,390.00 Q 637.32,393.03 643.20,390.00 Q 637.32,386.97 630.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,390.00 Q 633.03,397.32 639.33,399.33 Q 637.32,393.03 630.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,390.00 Q 626.97,397.32 630.00,403.20 Q 633.03,397.32 630.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,390.00 Q 622.68,393.03 620.67,399.33 Q 626.97,397.32 630.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,390.00 Q 622.68,386.97 616.80,390.00 Q 622.68,393.03 630.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,390.00 Q 626.97,382.68 620.67,380.67 Q 622.68,386.97 630.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,390.00 Q 633.03,382.68 630.00,376.80 Q 626.97,382.68 630.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,390.00 Q 637.32,386.97 639.33,380.67 Q 633.03,382.68 630.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,390.00 Q 630.93,393.48 635.09,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,390.00 Q 626.52,390.93 624.91,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,390.00 Q 629.07,386.52 624.91,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,390.00 Q 633.48,389.07 635.09,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="630.0" cy="390.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 630.00,405.12 C 623.60,398.72 616.74,391.86 614.88,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,374.88 C 636.40,381.28 643.26,388.14 645.12,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 664.80,390.00 C 675.78,379.02 686.58,368.22 690.00,364.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 715.20,390.00 C 704.22,400.98 693.42,411.78 690.00,415.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 690.00,390.00 Q 697.32,393.03 703.20,390.00 Q 697.32,386.97 690.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,390.00 Q 693.03,397.32 699.33,399.33 Q 697.32,393.03 690.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,390.00 Q 686.97,397.32 690.00,403.20 Q 693.03,397.32 690.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,390.00 Q 682.68,393.03 680.67,399.33 Q 686.97,397.32 690.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,390.00 Q 682.68,386.97 676.80,390.00 Q 682.68,393.03 690.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,390.00 Q 686.97,382.68 680.67,380.67 Q 682.68,386.97 690.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,390.00 Q 693.03,382.68 690.00,376.80 Q 686.97,382.68 690.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,390.00 Q 697.32,386.97 699.33,380.67 Q 693.03,382.68 690.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,390.00 Q 690.93,393.48 695.09,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,390.00 Q 686.52,390.93 684.91,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,390.00 Q 689.07,386.52 684.91,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,390.00 Q 693.48,389.07 695.09,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="690.0" cy="390.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 690.00,374.88 C 696.40,381.28 703.26,388.14 705.12,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,405.12 C 683.60,398.72 676.74,391.86 674.88,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 750.00,415.20 C 739.02,404.22 728.22,393.42 724.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,364.80 C 760.98,375.78 771.78,386.58 775.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 734.88,390.00 C 741.28,383.60 748.14,376.74 750.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 765.12,390.00 C 758.72,396.40 751.86,403.26 750.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 810.00,415.20 C 799.02,404.22 788.22,393.42 784.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,364.80 C 820.98,375.78 831.78,386.58 835.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 810.00,390.00 Q 817.32,393.03 823.20,390.00 Q 817.32,386.97 810.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,390.00 Q 813.03,397.32 819.33,399.33 Q 817.32,393.03 810.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,390.00 Q 806.97,397.32 810.00,403.20 Q 813.03,397.32 810.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,390.00 Q 802.68,393.03 800.67,399.33 Q 806.97,397.32 810.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,390.00 Q 802.68,386.97 796.80,390.00 Q 802.68,393.03 810.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,390.00 Q 806.97,382.68 800.67,380.67 Q 802.68,386.97 810.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,390.00 Q 813.03,382.68 810.00,376.80 Q 806.97,382.68 810.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,390.00 Q 817.32,386.97 819.33,380.67 Q 813.03,382.68 810.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,390.00 Q 810.93,393.48 815.09,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,390.00 Q 806.52,390.93 804.91,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,390.00 Q 809.07,386.52 804.91,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,390.00 Q 813.48,389.07 815.09,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="810.0" cy="390.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 794.88,390.00 C 801.28,383.60 808.14,376.74 810.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 825.12,390.00 C 818.72,396.40 811.86,403.26 810.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 870.00,364.80 C 880.98,375.78 891.78,386.58 895.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,415.20 C 859.02,404.22 848.22,393.42 844.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,390.00 Q 877.32,393.03 883.20,390.00 Q 877.32,386.97 870.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,390.00 Q 873.03,397.32 879.33,399.33 Q 877.32,393.03 870.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,390.00 Q 866.97,397.32 870.00,403.20 Q 873.03,397.32 870.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,390.00 Q 862.68,393.03 860.67,399.33 Q 866.97,397.32 870.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,390.00 Q 862.68,386.97 856.80,390.00 Q 862.68,393.03 870.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,390.00 Q 866.97,382.68 860.67,380.67 Q 862.68,386.97 870.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,390.00 Q 873.03,382.68 870.00,376.80 Q 866.97,382.68 870.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,390.00 Q 877.32,386.97 879.33,380.67 Q 873.03,382.68 870.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,390.00 Q 870.93,393.48 875.09,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,390.00 Q 866.52,390.93 864.91,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,390.00 Q 869.07,386.52 864.91,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,390.00 Q 873.48,389.07 875.09,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="390.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 885.12,390.00 C 878.72,396.40 871.86,403.26 870.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 854.88,390.00 C 861.28,383.60 868.14,376.74 870.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 904.80,390.00 C 915.78,379.02 926.58,368.22 930.00,364.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 955.20,390.00 C 944.22,400.98 933.42,411.78 930.00,415.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,390.00 Q 937.32,393.03 943.20,390.00 Q 937.32,386.97 930.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,390.00 Q 933.03,397.32 939.33,399.33 Q 937.32,393.03 930.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,390.00 Q 926.97,397.32 930.00,403.20 Q 933.03,397.32 930.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,390.00 Q 922.68,393.03 920.67,399.33 Q 926.97,397.32 930.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,390.00 Q 922.68,386.97 916.80,390.00 Q 922.68,393.03 930.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,390.00 Q 926.97,382.68 920.67,380.67 Q 922.68,386.97 930.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,390.00 Q 933.03,382.68 930.00,376.80 Q 926.97,382.68 930.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,390.00 Q 937.32,386.97 939.33,380.67 Q 933.03,382.68 930.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,390.00 Q 930.93,393.48 935.09,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,390.00 Q 926.52,390.93 924.91,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,390.00 Q 929.07,386.52 924.91,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,390.00 Q 933.48,389.07 935.09,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="390.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 930.00,374.88 C 936.40,381.28 943.26,388.14 945.12,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,405.12 C 923.60,398.72 916.74,391.86 914.88,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,364.80 C 1000.98,375.78 1011.78,386.58 1015.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,415.20 C 979.02,404.22 968.22,393.42 964.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1005.12,390.00 C 998.72,396.40 991.86,403.26 990.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 974.88,390.00 C 981.28,383.60 988.14,376.74 990.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1050.00,364.80 C 1060.98,375.78 1071.78,386.58 1075.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,415.20 C 1039.02,404.22 1028.22,393.42 1024.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1065.12,390.00 C 1058.72,396.40 1051.86,403.26 1050.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1034.88,390.00 C 1041.28,383.60 1048.14,376.74 1050.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1084.80,390.00 C 1095.78,379.02 1106.58,368.22 1110.00,364.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1135.20,390.00 C 1124.22,400.98 1113.42,411.78 1110.00,415.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1110.00,374.88 C 1116.40,381.28 1123.26,388.14 1125.12,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,405.12 C 1103.60,398.72 1096.74,391.86 1094.88,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1144.80,390.00 C 1155.78,379.02 1166.58,368.22 1170.00,364.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1195.20,390.00 C 1184.22,400.98 1173.42,411.78 1170.00,415.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1170.00,390.00 Q 1177.32,393.03 1183.20,390.00 Q 1177.32,386.97 1170.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,390.00 Q 1173.03,397.32 1179.33,399.33 Q 1177.32,393.03 1170.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,390.00 Q 1166.97,397.32 1170.00,403.20 Q 1173.03,397.32 1170.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,390.00 Q 1162.68,393.03 1160.67,399.33 Q 1166.97,397.32 1170.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,390.00 Q 1162.68,386.97 1156.80,390.00 Q 1162.68,393.03 1170.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,390.00 Q 1166.97,382.68 1160.67,380.67 Q 1162.68,386.97 1170.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,390.00 Q 1173.03,382.68 1170.00,376.80 Q 1166.97,382.68 1170.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,390.00 Q 1177.32,386.97 1179.33,380.67 Q 1173.03,382.68 1170.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,390.00 Q 1170.93,393.48 1175.09,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,390.00 Q 1166.52,390.93 1164.91,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,390.00 Q 1169.07,386.52 1164.91,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,390.00 Q 1173.48,389.07 1175.09,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1170.0" cy="390.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1170.00,374.88 C 1176.40,381.28 1183.26,388.14 1185.12,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,405.12 C 1163.60,398.72 1156.74,391.86 1154.88,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,415.20 C 1219.02,404.22 1208.22,393.42 1204.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,364.80 C 1240.98,375.78 1251.78,386.58 1255.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1214.88,390.00 C 1221.28,383.60 1228.14,376.74 1230.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1245.12,390.00 C 1238.72,396.40 1231.86,403.26 1230.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1290.00,415.20 C 1279.02,404.22 1268.22,393.42 1264.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,364.80 C 1300.98,375.78 1311.78,386.58 1315.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1274.88,390.00 C 1281.28,383.60 1288.14,376.74 1290.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1305.12,390.00 C 1298.72,396.40 1291.86,403.26 1290.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1350.00,364.80 C 1360.98,375.78 1371.78,386.58 1375.20,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,415.20 C 1339.02,404.22 1328.22,393.42 1324.80,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1350.00,390.00 Q 1357.32,393.03 1363.20,390.00 Q 1357.32,386.97 1350.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,390.00 Q 1353.03,397.32 1359.33,399.33 Q 1357.32,393.03 1350.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,390.00 Q 1346.97,397.32 1350.00,403.20 Q 1353.03,397.32 1350.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,390.00 Q 1342.68,393.03 1340.67,399.33 Q 1346.97,397.32 1350.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,390.00 Q 1342.68,386.97 1336.80,390.00 Q 1342.68,393.03 1350.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,390.00 Q 1346.97,382.68 1340.67,380.67 Q 1342.68,386.97 1350.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,390.00 Q 1353.03,382.68 1350.00,376.80 Q 1346.97,382.68 1350.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,390.00 Q 1357.32,386.97 1359.33,380.67 Q 1353.03,382.68 1350.00,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,390.00 Q 1350.93,393.48 1355.09,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,390.00 Q 1346.52,390.93 1344.91,395.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,390.00 Q 1349.07,386.52 1344.91,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,390.00 Q 1353.48,389.07 1355.09,384.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1350.0" cy="390.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1365.12,390.00 C 1358.72,396.40 1351.86,403.26 1350.00,405.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1334.88,390.00 C 1341.28,383.60 1348.14,376.74 1350.00,374.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,424.80 C 160.98,435.78 171.78,446.58 175.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,475.20 C 139.02,464.22 128.22,453.42 124.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,450.00 Q 157.32,453.03 163.20,450.00 Q 157.32,446.97 150.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,450.00 Q 153.03,457.32 159.33,459.33 Q 157.32,453.03 150.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,450.00 Q 146.97,457.32 150.00,463.20 Q 153.03,457.32 150.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,450.00 Q 142.68,453.03 140.67,459.33 Q 146.97,457.32 150.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,450.00 Q 142.68,446.97 136.80,450.00 Q 142.68,453.03 150.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,450.00 Q 146.97,442.68 140.67,440.67 Q 142.68,446.97 150.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,450.00 Q 153.03,442.68 150.00,436.80 Q 146.97,442.68 150.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,450.00 Q 157.32,446.97 159.33,440.67 Q 153.03,442.68 150.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,450.00 Q 150.93,453.48 155.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,450.00 Q 146.52,450.93 144.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,450.00 Q 149.07,446.52 144.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,450.00 Q 153.48,449.07 155.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 165.12,450.00 C 158.72,456.40 151.86,463.26 150.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 134.88,450.00 C 141.28,443.60 148.14,436.74 150.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 235.20,450.00 C 224.22,460.98 213.42,471.78 210.00,475.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 184.80,450.00 C 195.78,439.02 206.58,428.22 210.00,424.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,465.12 C 203.60,458.72 196.74,451.86 194.88,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,434.88 C 216.40,441.28 223.26,448.14 225.12,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,424.80 C 280.98,435.78 291.78,446.58 295.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,475.20 C 259.02,464.22 248.22,453.42 244.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 285.12,450.00 C 278.72,456.40 271.86,463.26 270.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 254.88,450.00 C 261.28,443.60 268.14,436.74 270.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,450.00 C 315.78,439.02 326.58,428.22 330.00,424.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,450.00 C 344.22,460.98 333.42,471.78 330.00,475.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 330.00,434.88 C 336.40,441.28 343.26,448.14 345.12,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,465.12 C 323.60,458.72 316.74,451.86 314.88,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,450.00 C 375.78,439.02 386.58,428.22 390.00,424.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,450.00 C 404.22,460.98 393.42,471.78 390.00,475.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 390.00,450.00 Q 397.32,453.03 403.20,450.00 Q 397.32,446.97 390.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,450.00 Q 393.03,457.32 399.33,459.33 Q 397.32,453.03 390.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,450.00 Q 386.97,457.32 390.00,463.20 Q 393.03,457.32 390.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,450.00 Q 382.68,453.03 380.67,459.33 Q 386.97,457.32 390.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,450.00 Q 382.68,446.97 376.80,450.00 Q 382.68,453.03 390.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,450.00 Q 386.97,442.68 380.67,440.67 Q 382.68,446.97 390.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,450.00 Q 393.03,442.68 390.00,436.80 Q 386.97,442.68 390.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,450.00 Q 397.32,446.97 399.33,440.67 Q 393.03,442.68 390.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,450.00 Q 390.93,453.48 395.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,450.00 Q 386.52,450.93 384.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,450.00 Q 389.07,446.52 384.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,450.00 Q 393.48,449.07 395.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="390.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 390.00,434.88 C 396.40,441.28 403.26,448.14 405.12,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,465.12 C 383.60,458.72 376.74,451.86 374.88,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 450.00,475.20 C 439.02,464.22 428.22,453.42 424.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,424.80 C 460.98,435.78 471.78,446.58 475.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 434.88,450.00 C 441.28,443.60 448.14,436.74 450.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 465.12,450.00 C 458.72,456.40 451.86,463.26 450.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,475.20 C 499.02,464.22 488.22,453.42 484.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,424.80 C 520.98,435.78 531.78,446.58 535.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,450.00 Q 517.32,453.03 523.20,450.00 Q 517.32,446.97 510.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,450.00 Q 513.03,457.32 519.33,459.33 Q 517.32,453.03 510.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,450.00 Q 506.97,457.32 510.00,463.20 Q 513.03,457.32 510.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,450.00 Q 502.68,453.03 500.67,459.33 Q 506.97,457.32 510.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,450.00 Q 502.68,446.97 496.80,450.00 Q 502.68,453.03 510.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,450.00 Q 506.97,442.68 500.67,440.67 Q 502.68,446.97 510.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,450.00 Q 513.03,442.68 510.00,436.80 Q 506.97,442.68 510.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,450.00 Q 517.32,446.97 519.33,440.67 Q 513.03,442.68 510.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,450.00 Q 510.93,453.48 515.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,450.00 Q 506.52,450.93 504.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,450.00 Q 509.07,446.52 504.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,450.00 Q 513.48,449.07 515.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 494.88,450.00 C 501.28,443.60 508.14,436.74 510.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 525.12,450.00 C 518.72,456.40 511.86,463.26 510.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 570.00,424.80 C 580.98,435.78 591.78,446.58 595.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,475.20 C 559.02,464.22 548.22,453.42 544.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 570.00,450.00 Q 577.32,453.03 583.20,450.00 Q 577.32,446.97 570.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,450.00 Q 573.03,457.32 579.33,459.33 Q 577.32,453.03 570.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,450.00 Q 566.97,457.32 570.00,463.20 Q 573.03,457.32 570.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,450.00 Q 562.68,453.03 560.67,459.33 Q 566.97,457.32 570.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,450.00 Q 562.68,446.97 556.80,450.00 Q 562.68,453.03 570.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,450.00 Q 566.97,442.68 560.67,440.67 Q 562.68,446.97 570.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,450.00 Q 573.03,442.68 570.00,436.80 Q 566.97,442.68 570.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,450.00 Q 577.32,446.97 579.33,440.67 Q 573.03,442.68 570.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,450.00 Q 570.93,453.48 575.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,450.00 Q 566.52,450.93 564.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,450.00 Q 569.07,446.52 564.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,450.00 Q 573.48,449.07 575.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="570.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 585.12,450.00 C 578.72,456.40 571.86,463.26 570.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 554.88,450.00 C 561.28,443.60 568.14,436.74 570.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,450.00 C 615.78,439.02 626.58,428.22 630.00,424.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,450.00 C 644.22,460.98 633.42,471.78 630.00,475.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 630.00,450.00 Q 637.32,453.03 643.20,450.00 Q 637.32,446.97 630.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,450.00 Q 633.03,457.32 639.33,459.33 Q 637.32,453.03 630.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,450.00 Q 626.97,457.32 630.00,463.20 Q 633.03,457.32 630.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,450.00 Q 622.68,453.03 620.67,459.33 Q 626.97,457.32 630.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,450.00 Q 622.68,446.97 616.80,450.00 Q 622.68,453.03 630.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,450.00 Q 626.97,442.68 620.67,440.67 Q 622.68,446.97 630.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,450.00 Q 633.03,442.68 630.00,436.80 Q 626.97,442.68 630.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,450.00 Q 637.32,446.97 639.33,440.67 Q 633.03,442.68 630.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,450.00 Q 630.93,453.48 635.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,450.00 Q 626.52,450.93 624.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,450.00 Q 629.07,446.52 624.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,450.00 Q 633.48,449.07 635.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="630.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 630.00,434.88 C 636.40,441.28 643.26,448.14 645.12,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,465.12 C 623.60,458.72 616.74,451.86 614.88,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 690.00,424.80 C 700.98,435.78 711.78,446.58 715.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,475.20 C 679.02,464.22 668.22,453.42 664.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 705.12,450.00 C 698.72,456.40 691.86,463.26 690.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 674.88,450.00 C 681.28,443.60 688.14,436.74 690.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 750.00,475.20 C 739.02,464.22 728.22,453.42 724.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,424.80 C 760.98,435.78 771.78,446.58 775.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 734.88,450.00 C 741.28,443.60 748.14,436.74 750.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 765.12,450.00 C 758.72,456.40 751.86,463.26 750.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 810.00,424.80 C 820.98,435.78 831.78,446.58 835.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,475.20 C 799.02,464.22 788.22,453.42 784.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 810.00,450.00 Q 817.32,453.03 823.20,450.00 Q 817.32,446.97 810.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,450.00 Q 813.03,457.32 819.33,459.33 Q 817.32,453.03 810.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,450.00 Q 806.97,457.32 810.00,463.20 Q 813.03,457.32 810.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,450.00 Q 802.68,453.03 800.67,459.33 Q 806.97,457.32 810.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,450.00 Q 802.68,446.97 796.80,450.00 Q 802.68,453.03 810.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,450.00 Q 806.97,442.68 800.67,440.67 Q 802.68,446.97 810.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,450.00 Q 813.03,442.68 810.00,436.80 Q 806.97,442.68 810.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,450.00 Q 817.32,446.97 819.33,440.67 Q 813.03,442.68 810.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,450.00 Q 810.93,453.48 815.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,450.00 Q 806.52,450.93 804.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,450.00 Q 809.07,446.52 804.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,450.00 Q 813.48,449.07 815.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="810.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 825.12,450.00 C 818.72,456.40 811.86,463.26 810.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 794.88,450.00 C 801.28,443.60 808.14,436.74 810.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 844.80,450.00 C 855.78,439.02 866.58,428.22 870.00,424.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 895.20,450.00 C 884.22,460.98 873.42,471.78 870.00,475.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,450.00 Q 877.32,453.03 883.20,450.00 Q 877.32,446.97 870.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,450.00 Q 873.03,457.32 879.33,459.33 Q 877.32,453.03 870.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,450.00 Q 866.97,457.32 870.00,463.20 Q 873.03,457.32 870.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,450.00 Q 862.68,453.03 860.67,459.33 Q 866.97,457.32 870.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,450.00 Q 862.68,446.97 856.80,450.00 Q 862.68,453.03 870.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,450.00 Q 866.97,442.68 860.67,440.67 Q 862.68,446.97 870.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,450.00 Q 873.03,442.68 870.00,436.80 Q 866.97,442.68 870.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,450.00 Q 877.32,446.97 879.33,440.67 Q 873.03,442.68 870.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,450.00 Q 870.93,453.48 875.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,450.00 Q 866.52,450.93 864.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,450.00 Q 869.07,446.52 864.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,450.00 Q 873.48,449.07 875.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 870.00,434.88 C 876.40,441.28 883.26,448.14 885.12,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,465.12 C 863.60,458.72 856.74,451.86 854.88,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 955.20,450.00 C 944.22,460.98 933.42,471.78 930.00,475.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 904.80,450.00 C 915.78,439.02 926.58,428.22 930.00,424.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,450.00 Q 937.32,453.03 943.20,450.00 Q 937.32,446.97 930.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,450.00 Q 933.03,457.32 939.33,459.33 Q 937.32,453.03 930.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,450.00 Q 926.97,457.32 930.00,463.20 Q 933.03,457.32 930.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,450.00 Q 922.68,453.03 920.67,459.33 Q 926.97,457.32 930.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,450.00 Q 922.68,446.97 916.80,450.00 Q 922.68,453.03 930.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,450.00 Q 926.97,442.68 920.67,440.67 Q 922.68,446.97 930.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,450.00 Q 933.03,442.68 930.00,436.80 Q 926.97,442.68 930.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,450.00 Q 937.32,446.97 939.33,440.67 Q 933.03,442.68 930.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,450.00 Q 930.93,453.48 935.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,450.00 Q 926.52,450.93 924.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,450.00 Q 929.07,446.52 924.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,450.00 Q 933.48,449.07 935.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 930.00,465.12 C 923.60,458.72 916.74,451.86 914.88,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,434.88 C 936.40,441.28 943.26,448.14 945.12,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,424.80 C 1000.98,435.78 1011.78,446.58 1015.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,475.20 C 979.02,464.22 968.22,453.42 964.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 990.00,450.00 Q 997.32,453.03 1003.20,450.00 Q 997.32,446.97 990.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,450.00 Q 993.03,457.32 999.33,459.33 Q 997.32,453.03 990.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,450.00 Q 986.97,457.32 990.00,463.20 Q 993.03,457.32 990.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,450.00 Q 982.68,453.03 980.67,459.33 Q 986.97,457.32 990.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,450.00 Q 982.68,446.97 976.80,450.00 Q 982.68,453.03 990.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,450.00 Q 986.97,442.68 980.67,440.67 Q 982.68,446.97 990.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,450.00 Q 993.03,442.68 990.00,436.80 Q 986.97,442.68 990.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,450.00 Q 997.32,446.97 999.33,440.67 Q 993.03,442.68 990.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,450.00 Q 990.93,453.48 995.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,450.00 Q 986.52,450.93 984.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,450.00 Q 989.07,446.52 984.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,450.00 Q 993.48,449.07 995.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="990.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1005.12,450.00 C 998.72,456.40 991.86,463.26 990.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 974.88,450.00 C 981.28,443.60 988.14,436.74 990.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1050.00,424.80 C 1060.98,435.78 1071.78,446.58 1075.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,475.20 C 1039.02,464.22 1028.22,453.42 1024.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1050.00,450.00 Q 1057.32,453.03 1063.20,450.00 Q 1057.32,446.97 1050.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,450.00 Q 1053.03,457.32 1059.33,459.33 Q 1057.32,453.03 1050.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,450.00 Q 1046.97,457.32 1050.00,463.20 Q 1053.03,457.32 1050.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,450.00 Q 1042.68,453.03 1040.67,459.33 Q 1046.97,457.32 1050.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,450.00 Q 1042.68,446.97 1036.80,450.00 Q 1042.68,453.03 1050.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,450.00 Q 1046.97,442.68 1040.67,440.67 Q 1042.68,446.97 1050.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,450.00 Q 1053.03,442.68 1050.00,436.80 Q 1046.97,442.68 1050.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,450.00 Q 1057.32,446.97 1059.33,440.67 Q 1053.03,442.68 1050.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,450.00 Q 1050.93,453.48 1055.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,450.00 Q 1046.52,450.93 1044.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,450.00 Q 1049.07,446.52 1044.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,450.00 Q 1053.48,449.07 1055.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1050.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1065.12,450.00 C 1058.72,456.40 1051.86,463.26 1050.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1034.88,450.00 C 1041.28,443.60 1048.14,436.74 1050.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1110.00,424.80 C 1120.98,435.78 1131.78,446.58 1135.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,475.20 C 1099.02,464.22 1088.22,453.42 1084.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1110.00,450.00 Q 1117.32,453.03 1123.20,450.00 Q 1117.32,446.97 1110.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,450.00 Q 1113.03,457.32 1119.33,459.33 Q 1117.32,453.03 1110.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,450.00 Q 1106.97,457.32 1110.00,463.20 Q 1113.03,457.32 1110.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,450.00 Q 1102.68,453.03 1100.67,459.33 Q 1106.97,457.32 1110.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,450.00 Q 1102.68,446.97 1096.80,450.00 Q 1102.68,453.03 1110.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,450.00 Q 1106.97,442.68 1100.67,440.67 Q 1102.68,446.97 1110.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,450.00 Q 1113.03,442.68 1110.00,436.80 Q 1106.97,442.68 1110.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,450.00 Q 1117.32,446.97 1119.33,440.67 Q 1113.03,442.68 1110.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,450.00 Q 1110.93,453.48 1115.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,450.00 Q 1106.52,450.93 1104.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,450.00 Q 1109.07,446.52 1104.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,450.00 Q 1113.48,449.07 1115.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1110.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1125.12,450.00 C 1118.72,456.40 1111.86,463.26 1110.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1094.88,450.00 C 1101.28,443.60 1108.14,436.74 1110.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1195.20,450.00 C 1184.22,460.98 1173.42,471.78 1170.00,475.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1144.80,450.00 C 1155.78,439.02 1166.58,428.22 1170.00,424.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1170.00,465.12 C 1163.60,458.72 1156.74,451.86 1154.88,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,434.88 C 1176.40,441.28 1183.26,448.14 1185.12,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,475.20 C 1219.02,464.22 1208.22,453.42 1204.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,424.80 C 1240.98,435.78 1251.78,446.58 1255.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1230.00,450.00 Q 1237.32,453.03 1243.20,450.00 Q 1237.32,446.97 1230.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,450.00 Q 1233.03,457.32 1239.33,459.33 Q 1237.32,453.03 1230.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,450.00 Q 1226.97,457.32 1230.00,463.20 Q 1233.03,457.32 1230.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,450.00 Q 1222.68,453.03 1220.67,459.33 Q 1226.97,457.32 1230.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,450.00 Q 1222.68,446.97 1216.80,450.00 Q 1222.68,453.03 1230.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,450.00 Q 1226.97,442.68 1220.67,440.67 Q 1222.68,446.97 1230.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,450.00 Q 1233.03,442.68 1230.00,436.80 Q 1226.97,442.68 1230.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,450.00 Q 1237.32,446.97 1239.33,440.67 Q 1233.03,442.68 1230.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,450.00 Q 1230.93,453.48 1235.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,450.00 Q 1226.52,450.93 1224.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,450.00 Q 1229.07,446.52 1224.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,450.00 Q 1233.48,449.07 1235.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1230.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1214.88,450.00 C 1221.28,443.60 1228.14,436.74 1230.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1245.12,450.00 C 1238.72,456.40 1231.86,463.26 1230.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1290.00,424.80 C 1300.98,435.78 1311.78,446.58 1315.20,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,475.20 C 1279.02,464.22 1268.22,453.42 1264.80,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1290.00,450.00 Q 1297.32,453.03 1303.20,450.00 Q 1297.32,446.97 1290.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,450.00 Q 1293.03,457.32 1299.33,459.33 Q 1297.32,453.03 1290.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,450.00 Q 1286.97,457.32 1290.00,463.20 Q 1293.03,457.32 1290.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,450.00 Q 1282.68,453.03 1280.67,459.33 Q 1286.97,457.32 1290.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,450.00 Q 1282.68,446.97 1276.80,450.00 Q 1282.68,453.03 1290.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,450.00 Q 1286.97,442.68 1280.67,440.67 Q 1282.68,446.97 1290.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,450.00 Q 1293.03,442.68 1290.00,436.80 Q 1286.97,442.68 1290.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,450.00 Q 1297.32,446.97 1299.33,440.67 Q 1293.03,442.68 1290.00,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,450.00 Q 1290.93,453.48 1295.09,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,450.00 Q 1286.52,450.93 1284.91,455.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,450.00 Q 1289.07,446.52 1284.91,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,450.00 Q 1293.48,449.07 1295.09,444.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1290.0" cy="450.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1305.12,450.00 C 1298.72,456.40 1291.86,463.26 1290.00,465.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1274.88,450.00 C 1281.28,443.60 1288.14,436.74 1290.00,434.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1324.80,450.00 C 1335.78,439.02 1346.58,428.22 1350.00,424.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1375.20,450.00 C 1364.22,460.98 1353.42,471.78 1350.00,475.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,434.88 C 1356.40,441.28 1363.26,448.14 1365.12,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,465.12 C 1343.60,458.72 1336.74,451.86 1334.88,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 175.20,510.00 C 164.22,520.98 153.42,531.78 150.00,535.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 124.80,510.00 C 135.78,499.02 146.58,488.22 150.00,484.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 150.00,525.12 C 143.60,518.72 136.74,511.86 134.88,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,494.88 C 156.40,501.28 163.26,508.14 165.12,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 184.80,510.00 C 195.78,499.02 206.58,488.22 210.00,484.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 235.20,510.00 C 224.22,520.98 213.42,531.78 210.00,535.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,494.88 C 216.40,501.28 223.26,508.14 225.12,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,525.12 C 203.60,518.72 196.74,511.86 194.88,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,484.80 C 280.98,495.78 291.78,506.58 295.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,535.20 C 259.02,524.22 248.22,513.42 244.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 270.00,510.00 Q 277.32,513.03 283.20,510.00 Q 277.32,506.97 270.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,510.00 Q 273.03,517.32 279.33,519.33 Q 277.32,513.03 270.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,510.00 Q 266.97,517.32 270.00,523.20 Q 273.03,517.32 270.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,510.00 Q 262.68,513.03 260.67,519.33 Q 266.97,517.32 270.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,510.00 Q 262.68,506.97 256.80,510.00 Q 262.68,513.03 270.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,510.00 Q 266.97,502.68 260.67,500.67 Q 262.68,506.97 270.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,510.00 Q 273.03,502.68 270.00,496.80 Q 266.97,502.68 270.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,510.00 Q 277.32,506.97 279.33,500.67 Q 273.03,502.68 270.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,510.00 Q 270.93,513.48 275.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,510.00 Q 266.52,510.93 264.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,510.00 Q 269.07,506.52 264.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,510.00 Q 273.48,509.07 275.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="270.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 285.12,510.00 C 278.72,516.40 271.86,523.26 270.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 254.88,510.00 C 261.28,503.60 268.14,496.74 270.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,510.00 C 315.78,499.02 326.58,488.22 330.00,484.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,510.00 C 344.22,520.98 333.42,531.78 330.00,535.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 330.00,510.00 Q 337.32,513.03 343.20,510.00 Q 337.32,506.97 330.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,510.00 Q 333.03,517.32 339.33,519.33 Q 337.32,513.03 330.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,510.00 Q 326.97,517.32 330.00,523.20 Q 333.03,517.32 330.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,510.00 Q 322.68,513.03 320.67,519.33 Q 326.97,517.32 330.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,510.00 Q 322.68,506.97 316.80,510.00 Q 322.68,513.03 330.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,510.00 Q 326.97,502.68 320.67,500.67 Q 322.68,506.97 330.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,510.00 Q 333.03,502.68 330.00,496.80 Q 326.97,502.68 330.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,510.00 Q 337.32,506.97 339.33,500.67 Q 333.03,502.68 330.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,510.00 Q 330.93,513.48 335.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,510.00 Q 326.52,510.93 324.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,510.00 Q 329.07,506.52 324.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,510.00 Q 333.48,509.07 335.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="330.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 330.00,494.88 C 336.40,501.28 343.26,508.14 345.12,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,525.12 C 323.60,518.72 316.74,511.86 314.88,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 390.00,484.80 C 400.98,495.78 411.78,506.58 415.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,535.20 C 379.02,524.22 368.22,513.42 364.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 405.12,510.00 C 398.72,516.40 391.86,523.26 390.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 374.88,510.00 C 381.28,503.60 388.14,496.74 390.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 450.00,535.20 C 439.02,524.22 428.22,513.42 424.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,484.80 C 460.98,495.78 471.78,506.58 475.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 450.00,510.00 Q 457.32,513.03 463.20,510.00 Q 457.32,506.97 450.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,510.00 Q 453.03,517.32 459.33,519.33 Q 457.32,513.03 450.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,510.00 Q 446.97,517.32 450.00,523.20 Q 453.03,517.32 450.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,510.00 Q 442.68,513.03 440.67,519.33 Q 446.97,517.32 450.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,510.00 Q 442.68,506.97 436.80,510.00 Q 442.68,513.03 450.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,510.00 Q 446.97,502.68 440.67,500.67 Q 442.68,506.97 450.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,510.00 Q 453.03,502.68 450.00,496.80 Q 446.97,502.68 450.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,510.00 Q 457.32,506.97 459.33,500.67 Q 453.03,502.68 450.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,510.00 Q 450.93,513.48 455.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,510.00 Q 446.52,510.93 444.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,510.00 Q 449.07,506.52 444.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,510.00 Q 453.48,509.07 455.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="450.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 434.88,510.00 C 441.28,503.60 448.14,496.74 450.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 465.12,510.00 C 458.72,516.40 451.86,523.26 450.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,484.80 C 520.98,495.78 531.78,506.58 535.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,535.20 C 499.02,524.22 488.22,513.42 484.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,510.00 Q 517.32,513.03 523.20,510.00 Q 517.32,506.97 510.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,510.00 Q 513.03,517.32 519.33,519.33 Q 517.32,513.03 510.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,510.00 Q 506.97,517.32 510.00,523.20 Q 513.03,517.32 510.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,510.00 Q 502.68,513.03 500.67,519.33 Q 506.97,517.32 510.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,510.00 Q 502.68,506.97 496.80,510.00 Q 502.68,513.03 510.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,510.00 Q 506.97,502.68 500.67,500.67 Q 502.68,506.97 510.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,510.00 Q 513.03,502.68 510.00,496.80 Q 506.97,502.68 510.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,510.00 Q 517.32,506.97 519.33,500.67 Q 513.03,502.68 510.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,510.00 Q 510.93,513.48 515.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,510.00 Q 506.52,510.93 504.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,510.00 Q 509.07,506.52 504.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,510.00 Q 513.48,509.07 515.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 525.12,510.00 C 518.72,516.40 511.86,523.26 510.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 494.88,510.00 C 501.28,503.60 508.14,496.74 510.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 595.20,510.00 C 584.22,520.98 573.42,531.78 570.00,535.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 544.80,510.00 C 555.78,499.02 566.58,488.22 570.00,484.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 570.00,510.00 Q 577.32,513.03 583.20,510.00 Q 577.32,506.97 570.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,510.00 Q 573.03,517.32 579.33,519.33 Q 577.32,513.03 570.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,510.00 Q 566.97,517.32 570.00,523.20 Q 573.03,517.32 570.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,510.00 Q 562.68,513.03 560.67,519.33 Q 566.97,517.32 570.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,510.00 Q 562.68,506.97 556.80,510.00 Q 562.68,513.03 570.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,510.00 Q 566.97,502.68 560.67,500.67 Q 562.68,506.97 570.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,510.00 Q 573.03,502.68 570.00,496.80 Q 566.97,502.68 570.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,510.00 Q 577.32,506.97 579.33,500.67 Q 573.03,502.68 570.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,510.00 Q 570.93,513.48 575.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,510.00 Q 566.52,510.93 564.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,510.00 Q 569.07,506.52 564.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,510.00 Q 573.48,509.07 575.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="570.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 570.00,525.12 C 563.60,518.72 556.74,511.86 554.88,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,494.88 C 576.40,501.28 583.26,508.14 585.12,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 630.00,535.20 C 619.02,524.22 608.22,513.42 604.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,484.80 C 640.98,495.78 651.78,506.58 655.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 614.88,510.00 C 621.28,503.60 628.14,496.74 630.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 645.12,510.00 C 638.72,516.40 631.86,523.26 630.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 690.00,535.20 C 679.02,524.22 668.22,513.42 664.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,484.80 C 700.98,495.78 711.78,506.58 715.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 674.88,510.00 C 681.28,503.60 688.14,496.74 690.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 705.12,510.00 C 698.72,516.40 691.86,523.26 690.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 750.00,484.80 C 760.98,495.78 771.78,506.58 775.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,535.20 C 739.02,524.22 728.22,513.42 724.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 750.00,510.00 Q 757.32,513.03 763.20,510.00 Q 757.32,506.97 750.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,510.00 Q 753.03,517.32 759.33,519.33 Q 757.32,513.03 750.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,510.00 Q 746.97,517.32 750.00,523.20 Q 753.03,517.32 750.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,510.00 Q 742.68,513.03 740.67,519.33 Q 746.97,517.32 750.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,510.00 Q 742.68,506.97 736.80,510.00 Q 742.68,513.03 750.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,510.00 Q 746.97,502.68 740.67,500.67 Q 742.68,506.97 750.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,510.00 Q 753.03,502.68 750.00,496.80 Q 746.97,502.68 750.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,510.00 Q 757.32,506.97 759.33,500.67 Q 753.03,502.68 750.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,510.00 Q 750.93,513.48 755.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,510.00 Q 746.52,510.93 744.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,510.00 Q 749.07,506.52 744.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,510.00 Q 753.48,509.07 755.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="750.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 765.12,510.00 C 758.72,516.40 751.86,523.26 750.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 734.88,510.00 C 741.28,503.60 748.14,496.74 750.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 810.00,484.80 C 820.98,495.78 831.78,506.58 835.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,535.20 C 799.02,524.22 788.22,513.42 784.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 825.12,510.00 C 818.72,516.40 811.86,523.26 810.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 794.88,510.00 C 801.28,503.60 808.14,496.74 810.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 870.00,535.20 C 859.02,524.22 848.22,513.42 844.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,484.80 C 880.98,495.78 891.78,506.58 895.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 854.88,510.00 C 861.28,503.60 868.14,496.74 870.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 885.12,510.00 C 878.72,516.40 871.86,523.26 870.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 930.00,535.20 C 919.02,524.22 908.22,513.42 904.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,484.80 C 940.98,495.78 951.78,506.58 955.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 914.88,510.00 C 921.28,503.60 928.14,496.74 930.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 945.12,510.00 C 938.72,516.40 931.86,523.26 930.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,535.20 C 979.02,524.22 968.22,513.42 964.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,484.80 C 1000.98,495.78 1011.78,506.58 1015.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 990.00,510.00 Q 997.32,513.03 1003.20,510.00 Q 997.32,506.97 990.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,510.00 Q 993.03,517.32 999.33,519.33 Q 997.32,513.03 990.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,510.00 Q 986.97,517.32 990.00,523.20 Q 993.03,517.32 990.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,510.00 Q 982.68,513.03 980.67,519.33 Q 986.97,517.32 990.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,510.00 Q 982.68,506.97 976.80,510.00 Q 982.68,513.03 990.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,510.00 Q 986.97,502.68 980.67,500.67 Q 982.68,506.97 990.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,510.00 Q 993.03,502.68 990.00,496.80 Q 986.97,502.68 990.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,510.00 Q 997.32,506.97 999.33,500.67 Q 993.03,502.68 990.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,510.00 Q 990.93,513.48 995.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,510.00 Q 986.52,510.93 984.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,510.00 Q 989.07,506.52 984.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,510.00 Q 993.48,509.07 995.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="990.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 974.88,510.00 C 981.28,503.60 988.14,496.74 990.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1005.12,510.00 C 998.72,516.40 991.86,523.26 990.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,510.00 C 1035.78,499.02 1046.58,488.22 1050.00,484.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,510.00 C 1064.22,520.98 1053.42,531.78 1050.00,535.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1050.00,510.00 Q 1057.32,513.03 1063.20,510.00 Q 1057.32,506.97 1050.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,510.00 Q 1053.03,517.32 1059.33,519.33 Q 1057.32,513.03 1050.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,510.00 Q 1046.97,517.32 1050.00,523.20 Q 1053.03,517.32 1050.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,510.00 Q 1042.68,513.03 1040.67,519.33 Q 1046.97,517.32 1050.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,510.00 Q 1042.68,506.97 1036.80,510.00 Q 1042.68,513.03 1050.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,510.00 Q 1046.97,502.68 1040.67,500.67 Q 1042.68,506.97 1050.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,510.00 Q 1053.03,502.68 1050.00,496.80 Q 1046.97,502.68 1050.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,510.00 Q 1057.32,506.97 1059.33,500.67 Q 1053.03,502.68 1050.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,510.00 Q 1050.93,513.48 1055.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,510.00 Q 1046.52,510.93 1044.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,510.00 Q 1049.07,506.52 1044.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,510.00 Q 1053.48,509.07 1055.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1050.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1050.00,494.88 C 1056.40,501.28 1063.26,508.14 1065.12,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,525.12 C 1043.60,518.72 1036.74,511.86 1034.88,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1110.00,535.20 C 1099.02,524.22 1088.22,513.42 1084.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,484.80 C 1120.98,495.78 1131.78,506.58 1135.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1094.88,510.00 C 1101.28,503.60 1108.14,496.74 1110.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1125.12,510.00 C 1118.72,516.40 1111.86,523.26 1110.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1170.00,535.20 C 1159.02,524.22 1148.22,513.42 1144.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,484.80 C 1180.98,495.78 1191.78,506.58 1195.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1170.00,510.00 Q 1177.32,513.03 1183.20,510.00 Q 1177.32,506.97 1170.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,510.00 Q 1173.03,517.32 1179.33,519.33 Q 1177.32,513.03 1170.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,510.00 Q 1166.97,517.32 1170.00,523.20 Q 1173.03,517.32 1170.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,510.00 Q 1162.68,513.03 1160.67,519.33 Q 1166.97,517.32 1170.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,510.00 Q 1162.68,506.97 1156.80,510.00 Q 1162.68,513.03 1170.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,510.00 Q 1166.97,502.68 1160.67,500.67 Q 1162.68,506.97 1170.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,510.00 Q 1173.03,502.68 1170.00,496.80 Q 1166.97,502.68 1170.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,510.00 Q 1177.32,506.97 1179.33,500.67 Q 1173.03,502.68 1170.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,510.00 Q 1170.93,513.48 1175.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,510.00 Q 1166.52,510.93 1164.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,510.00 Q 1169.07,506.52 1164.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,510.00 Q 1173.48,509.07 1175.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1170.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1154.88,510.00 C 1161.28,503.60 1168.14,496.74 1170.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1185.12,510.00 C 1178.72,516.40 1171.86,523.26 1170.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,484.80 C 1240.98,495.78 1251.78,506.58 1255.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,535.20 C 1219.02,524.22 1208.22,513.42 1204.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1230.00,510.00 Q 1237.32,513.03 1243.20,510.00 Q 1237.32,506.97 1230.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,510.00 Q 1233.03,517.32 1239.33,519.33 Q 1237.32,513.03 1230.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,510.00 Q 1226.97,517.32 1230.00,523.20 Q 1233.03,517.32 1230.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,510.00 Q 1222.68,513.03 1220.67,519.33 Q 1226.97,517.32 1230.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,510.00 Q 1222.68,506.97 1216.80,510.00 Q 1222.68,513.03 1230.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,510.00 Q 1226.97,502.68 1220.67,500.67 Q 1222.68,506.97 1230.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,510.00 Q 1233.03,502.68 1230.00,496.80 Q 1226.97,502.68 1230.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,510.00 Q 1237.32,506.97 1239.33,500.67 Q 1233.03,502.68 1230.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,510.00 Q 1230.93,513.48 1235.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,510.00 Q 1226.52,510.93 1224.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,510.00 Q 1229.07,506.52 1224.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,510.00 Q 1233.48,509.07 1235.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1230.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1245.12,510.00 C 1238.72,516.40 1231.86,523.26 1230.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1214.88,510.00 C 1221.28,503.60 1228.14,496.74 1230.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1264.80,510.00 C 1275.78,499.02 1286.58,488.22 1290.00,484.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1315.20,510.00 C 1304.22,520.98 1293.42,531.78 1290.00,535.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1290.00,510.00 Q 1297.32,513.03 1303.20,510.00 Q 1297.32,506.97 1290.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,510.00 Q 1293.03,517.32 1299.33,519.33 Q 1297.32,513.03 1290.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,510.00 Q 1286.97,517.32 1290.00,523.20 Q 1293.03,517.32 1290.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,510.00 Q 1282.68,513.03 1280.67,519.33 Q 1286.97,517.32 1290.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,510.00 Q 1282.68,506.97 1276.80,510.00 Q 1282.68,513.03 1290.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,510.00 Q 1286.97,502.68 1280.67,500.67 Q 1282.68,506.97 1290.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,510.00 Q 1293.03,502.68 1290.00,496.80 Q 1286.97,502.68 1290.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,510.00 Q 1297.32,506.97 1299.33,500.67 Q 1293.03,502.68 1290.00,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,510.00 Q 1290.93,513.48 1295.09,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,510.00 Q 1286.52,510.93 1284.91,515.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,510.00 Q 1289.07,506.52 1284.91,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,510.00 Q 1293.48,509.07 1295.09,504.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1290.0" cy="510.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1290.00,494.88 C 1296.40,501.28 1303.26,508.14 1305.12,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,525.12 C 1283.60,518.72 1276.74,511.86 1274.88,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1350.00,484.80 C 1360.98,495.78 1371.78,506.58 1375.20,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,535.20 C 1339.02,524.22 1328.22,513.42 1324.80,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1365.12,510.00 C 1358.72,516.40 1351.86,523.26 1350.00,525.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1334.88,510.00 C 1341.28,503.60 1348.14,496.74 1350.00,494.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,595.20 C 139.02,584.22 128.22,573.42 124.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,544.80 C 160.98,555.78 171.78,566.58 175.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,570.00 Q 157.32,573.03 163.20,570.00 Q 157.32,566.97 150.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,570.00 Q 153.03,577.32 159.33,579.33 Q 157.32,573.03 150.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,570.00 Q 146.97,577.32 150.00,583.20 Q 153.03,577.32 150.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,570.00 Q 142.68,573.03 140.67,579.33 Q 146.97,577.32 150.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,570.00 Q 142.68,566.97 136.80,570.00 Q 142.68,573.03 150.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,570.00 Q 146.97,562.68 140.67,560.67 Q 142.68,566.97 150.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,570.00 Q 153.03,562.68 150.00,556.80 Q 146.97,562.68 150.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,570.00 Q 157.32,566.97 159.33,560.67 Q 153.03,562.68 150.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,570.00 Q 150.93,573.48 155.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,570.00 Q 146.52,570.93 144.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,570.00 Q 149.07,566.52 144.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,570.00 Q 153.48,569.07 155.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 134.88,570.00 C 141.28,563.60 148.14,556.74 150.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 165.12,570.00 C 158.72,576.40 151.86,583.26 150.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 210.00,544.80 C 220.98,555.78 231.78,566.58 235.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,595.20 C 199.02,584.22 188.22,573.42 184.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 210.00,570.00 Q 217.32,573.03 223.20,570.00 Q 217.32,566.97 210.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,570.00 Q 213.03,577.32 219.33,579.33 Q 217.32,573.03 210.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,570.00 Q 206.97,577.32 210.00,583.20 Q 213.03,577.32 210.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,570.00 Q 202.68,573.03 200.67,579.33 Q 206.97,577.32 210.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,570.00 Q 202.68,566.97 196.80,570.00 Q 202.68,573.03 210.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,570.00 Q 206.97,562.68 200.67,560.67 Q 202.68,566.97 210.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,570.00 Q 213.03,562.68 210.00,556.80 Q 206.97,562.68 210.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,570.00 Q 217.32,566.97 219.33,560.67 Q 213.03,562.68 210.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,570.00 Q 210.93,573.48 215.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,570.00 Q 206.52,570.93 204.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,570.00 Q 209.07,566.52 204.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,570.00 Q 213.48,569.07 215.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="210.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 225.12,570.00 C 218.72,576.40 211.86,583.26 210.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 194.88,570.00 C 201.28,563.60 208.14,556.74 210.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 244.80,570.00 C 255.78,559.02 266.58,548.22 270.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 295.20,570.00 C 284.22,580.98 273.42,591.78 270.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 270.00,570.00 Q 277.32,573.03 283.20,570.00 Q 277.32,566.97 270.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,570.00 Q 273.03,577.32 279.33,579.33 Q 277.32,573.03 270.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,570.00 Q 266.97,577.32 270.00,583.20 Q 273.03,577.32 270.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,570.00 Q 262.68,573.03 260.67,579.33 Q 266.97,577.32 270.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,570.00 Q 262.68,566.97 256.80,570.00 Q 262.68,573.03 270.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,570.00 Q 266.97,562.68 260.67,560.67 Q 262.68,566.97 270.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,570.00 Q 273.03,562.68 270.00,556.80 Q 266.97,562.68 270.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,570.00 Q 277.32,566.97 279.33,560.67 Q 273.03,562.68 270.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,570.00 Q 270.93,573.48 275.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,570.00 Q 266.52,570.93 264.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,570.00 Q 269.07,566.52 264.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,570.00 Q 273.48,569.07 275.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="270.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 270.00,554.88 C 276.40,561.28 283.26,568.14 285.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,585.12 C 263.60,578.72 256.74,571.86 254.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 355.20,570.00 C 344.22,580.98 333.42,591.78 330.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 304.80,570.00 C 315.78,559.02 326.58,548.22 330.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 330.00,570.00 Q 337.32,573.03 343.20,570.00 Q 337.32,566.97 330.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,570.00 Q 333.03,577.32 339.33,579.33 Q 337.32,573.03 330.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,570.00 Q 326.97,577.32 330.00,583.20 Q 333.03,577.32 330.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,570.00 Q 322.68,573.03 320.67,579.33 Q 326.97,577.32 330.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,570.00 Q 322.68,566.97 316.80,570.00 Q 322.68,573.03 330.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,570.00 Q 326.97,562.68 320.67,560.67 Q 322.68,566.97 330.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,570.00 Q 333.03,562.68 330.00,556.80 Q 326.97,562.68 330.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,570.00 Q 337.32,566.97 339.33,560.67 Q 333.03,562.68 330.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,570.00 Q 330.93,573.48 335.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,570.00 Q 326.52,570.93 324.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,570.00 Q 329.07,566.52 324.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,570.00 Q 333.48,569.07 335.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="330.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 330.00,585.12 C 323.60,578.72 316.74,571.86 314.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,554.88 C 336.40,561.28 343.26,568.14 345.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 390.00,544.80 C 400.98,555.78 411.78,566.58 415.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,595.20 C 379.02,584.22 368.22,573.42 364.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 390.00,570.00 Q 397.32,573.03 403.20,570.00 Q 397.32,566.97 390.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,570.00 Q 393.03,577.32 399.33,579.33 Q 397.32,573.03 390.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,570.00 Q 386.97,577.32 390.00,583.20 Q 393.03,577.32 390.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,570.00 Q 382.68,573.03 380.67,579.33 Q 386.97,577.32 390.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,570.00 Q 382.68,566.97 376.80,570.00 Q 382.68,573.03 390.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,570.00 Q 386.97,562.68 380.67,560.67 Q 382.68,566.97 390.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,570.00 Q 393.03,562.68 390.00,556.80 Q 386.97,562.68 390.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,570.00 Q 397.32,566.97 399.33,560.67 Q 393.03,562.68 390.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,570.00 Q 390.93,573.48 395.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,570.00 Q 386.52,570.93 384.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,570.00 Q 389.07,566.52 384.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,570.00 Q 393.48,569.07 395.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="390.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 405.12,570.00 C 398.72,576.40 391.86,583.26 390.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 374.88,570.00 C 381.28,563.60 388.14,556.74 390.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 450.00,544.80 C 460.98,555.78 471.78,566.58 475.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,595.20 C 439.02,584.22 428.22,573.42 424.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 450.00,570.00 Q 457.32,573.03 463.20,570.00 Q 457.32,566.97 450.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,570.00 Q 453.03,577.32 459.33,579.33 Q 457.32,573.03 450.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,570.00 Q 446.97,577.32 450.00,583.20 Q 453.03,577.32 450.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,570.00 Q 442.68,573.03 440.67,579.33 Q 446.97,577.32 450.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,570.00 Q 442.68,566.97 436.80,570.00 Q 442.68,573.03 450.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,570.00 Q 446.97,562.68 440.67,560.67 Q 442.68,566.97 450.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,570.00 Q 453.03,562.68 450.00,556.80 Q 446.97,562.68 450.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,570.00 Q 457.32,566.97 459.33,560.67 Q 453.03,562.68 450.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,570.00 Q 450.93,573.48 455.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,570.00 Q 446.52,570.93 444.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,570.00 Q 449.07,566.52 444.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,570.00 Q 453.48,569.07 455.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="450.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 465.12,570.00 C 458.72,576.40 451.86,583.26 450.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 434.88,570.00 C 441.28,563.60 448.14,556.74 450.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,544.80 C 520.98,555.78 531.78,566.58 535.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,595.20 C 499.02,584.22 488.22,573.42 484.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,570.00 Q 517.32,573.03 523.20,570.00 Q 517.32,566.97 510.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,570.00 Q 513.03,577.32 519.33,579.33 Q 517.32,573.03 510.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,570.00 Q 506.97,577.32 510.00,583.20 Q 513.03,577.32 510.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,570.00 Q 502.68,573.03 500.67,579.33 Q 506.97,577.32 510.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,570.00 Q 502.68,566.97 496.80,570.00 Q 502.68,573.03 510.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,570.00 Q 506.97,562.68 500.67,560.67 Q 502.68,566.97 510.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,570.00 Q 513.03,562.68 510.00,556.80 Q 506.97,562.68 510.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,570.00 Q 517.32,566.97 519.33,560.67 Q 513.03,562.68 510.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,570.00 Q 510.93,573.48 515.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,570.00 Q 506.52,570.93 504.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,570.00 Q 509.07,566.52 504.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,570.00 Q 513.48,569.07 515.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 525.12,570.00 C 518.72,576.40 511.86,583.26 510.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 494.88,570.00 C 501.28,563.60 508.14,556.74 510.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 595.20,570.00 C 584.22,580.98 573.42,591.78 570.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 544.80,570.00 C 555.78,559.02 566.58,548.22 570.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 570.00,585.12 C 563.60,578.72 556.74,571.86 554.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,554.88 C 576.40,561.28 583.26,568.14 585.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 630.00,595.20 C 619.02,584.22 608.22,573.42 604.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,544.80 C 640.98,555.78 651.78,566.58 655.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 630.00,570.00 Q 637.32,573.03 643.20,570.00 Q 637.32,566.97 630.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,570.00 Q 633.03,577.32 639.33,579.33 Q 637.32,573.03 630.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,570.00 Q 626.97,577.32 630.00,583.20 Q 633.03,577.32 630.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,570.00 Q 622.68,573.03 620.67,579.33 Q 626.97,577.32 630.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,570.00 Q 622.68,566.97 616.80,570.00 Q 622.68,573.03 630.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,570.00 Q 626.97,562.68 620.67,560.67 Q 622.68,566.97 630.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,570.00 Q 633.03,562.68 630.00,556.80 Q 626.97,562.68 630.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,570.00 Q 637.32,566.97 639.33,560.67 Q 633.03,562.68 630.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,570.00 Q 630.93,573.48 635.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,570.00 Q 626.52,570.93 624.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,570.00 Q 629.07,566.52 624.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,570.00 Q 633.48,569.07 635.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="630.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 614.88,570.00 C 621.28,563.60 628.14,556.74 630.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 645.12,570.00 C 638.72,576.40 631.86,583.26 630.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 690.00,544.80 C 700.98,555.78 711.78,566.58 715.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,595.20 C 679.02,584.22 668.22,573.42 664.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 690.00,570.00 Q 697.32,573.03 703.20,570.00 Q 697.32,566.97 690.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,570.00 Q 693.03,577.32 699.33,579.33 Q 697.32,573.03 690.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,570.00 Q 686.97,577.32 690.00,583.20 Q 693.03,577.32 690.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,570.00 Q 682.68,573.03 680.67,579.33 Q 686.97,577.32 690.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,570.00 Q 682.68,566.97 676.80,570.00 Q 682.68,573.03 690.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,570.00 Q 686.97,562.68 680.67,560.67 Q 682.68,566.97 690.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,570.00 Q 693.03,562.68 690.00,556.80 Q 686.97,562.68 690.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,570.00 Q 697.32,566.97 699.33,560.67 Q 693.03,562.68 690.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,570.00 Q 690.93,573.48 695.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,570.00 Q 686.52,570.93 684.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,570.00 Q 689.07,566.52 684.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,570.00 Q 693.48,569.07 695.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="690.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 705.12,570.00 C 698.72,576.40 691.86,583.26 690.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 674.88,570.00 C 681.28,563.60 688.14,556.74 690.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 775.20,570.00 C 764.22,580.98 753.42,591.78 750.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 724.80,570.00 C 735.78,559.02 746.58,548.22 750.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 750.00,570.00 Q 757.32,573.03 763.20,570.00 Q 757.32,566.97 750.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,570.00 Q 753.03,577.32 759.33,579.33 Q 757.32,573.03 750.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,570.00 Q 746.97,577.32 750.00,583.20 Q 753.03,577.32 750.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,570.00 Q 742.68,573.03 740.67,579.33 Q 746.97,577.32 750.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,570.00 Q 742.68,566.97 736.80,570.00 Q 742.68,573.03 750.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,570.00 Q 746.97,562.68 740.67,560.67 Q 742.68,566.97 750.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,570.00 Q 753.03,562.68 750.00,556.80 Q 746.97,562.68 750.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,570.00 Q 757.32,566.97 759.33,560.67 Q 753.03,562.68 750.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,570.00 Q 750.93,573.48 755.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,570.00 Q 746.52,570.93 744.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,570.00 Q 749.07,566.52 744.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,570.00 Q 753.48,569.07 755.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="750.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 750.00,585.12 C 743.60,578.72 736.74,571.86 734.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,554.88 C 756.40,561.28 763.26,568.14 765.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 835.20,570.00 C 824.22,580.98 813.42,591.78 810.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 784.80,570.00 C 795.78,559.02 806.58,548.22 810.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 810.00,570.00 Q 817.32,573.03 823.20,570.00 Q 817.32,566.97 810.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,570.00 Q 813.03,577.32 819.33,579.33 Q 817.32,573.03 810.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,570.00 Q 806.97,577.32 810.00,583.20 Q 813.03,577.32 810.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,570.00 Q 802.68,573.03 800.67,579.33 Q 806.97,577.32 810.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,570.00 Q 802.68,566.97 796.80,570.00 Q 802.68,573.03 810.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,570.00 Q 806.97,562.68 800.67,560.67 Q 802.68,566.97 810.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,570.00 Q 813.03,562.68 810.00,556.80 Q 806.97,562.68 810.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,570.00 Q 817.32,566.97 819.33,560.67 Q 813.03,562.68 810.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,570.00 Q 810.93,573.48 815.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,570.00 Q 806.52,570.93 804.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,570.00 Q 809.07,566.52 804.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,570.00 Q 813.48,569.07 815.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="810.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 810.00,585.12 C 803.60,578.72 796.74,571.86 794.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,554.88 C 816.40,561.28 823.26,568.14 825.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 870.00,544.80 C 880.98,555.78 891.78,566.58 895.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,595.20 C 859.02,584.22 848.22,573.42 844.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,570.00 Q 877.32,573.03 883.20,570.00 Q 877.32,566.97 870.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,570.00 Q 873.03,577.32 879.33,579.33 Q 877.32,573.03 870.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,570.00 Q 866.97,577.32 870.00,583.20 Q 873.03,577.32 870.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,570.00 Q 862.68,573.03 860.67,579.33 Q 866.97,577.32 870.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,570.00 Q 862.68,566.97 856.80,570.00 Q 862.68,573.03 870.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,570.00 Q 866.97,562.68 860.67,560.67 Q 862.68,566.97 870.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,570.00 Q 873.03,562.68 870.00,556.80 Q 866.97,562.68 870.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,570.00 Q 877.32,566.97 879.33,560.67 Q 873.03,562.68 870.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,570.00 Q 870.93,573.48 875.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,570.00 Q 866.52,570.93 864.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,570.00 Q 869.07,566.52 864.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,570.00 Q 873.48,569.07 875.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 885.12,570.00 C 878.72,576.40 871.86,583.26 870.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 854.88,570.00 C 861.28,563.60 868.14,556.74 870.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 930.00,544.80 C 940.98,555.78 951.78,566.58 955.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,595.20 C 919.02,584.22 908.22,573.42 904.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,570.00 Q 937.32,573.03 943.20,570.00 Q 937.32,566.97 930.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,570.00 Q 933.03,577.32 939.33,579.33 Q 937.32,573.03 930.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,570.00 Q 926.97,577.32 930.00,583.20 Q 933.03,577.32 930.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,570.00 Q 922.68,573.03 920.67,579.33 Q 926.97,577.32 930.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,570.00 Q 922.68,566.97 916.80,570.00 Q 922.68,573.03 930.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,570.00 Q 926.97,562.68 920.67,560.67 Q 922.68,566.97 930.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,570.00 Q 933.03,562.68 930.00,556.80 Q 926.97,562.68 930.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,570.00 Q 937.32,566.97 939.33,560.67 Q 933.03,562.68 930.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,570.00 Q 930.93,573.48 935.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,570.00 Q 926.52,570.93 924.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,570.00 Q 929.07,566.52 924.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,570.00 Q 933.48,569.07 935.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 945.12,570.00 C 938.72,576.40 931.86,583.26 930.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 914.88,570.00 C 921.28,563.60 928.14,556.74 930.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 964.80,570.00 C 975.78,559.02 986.58,548.22 990.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1015.20,570.00 C 1004.22,580.98 993.42,591.78 990.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 990.00,554.88 C 996.40,561.28 1003.26,568.14 1005.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,585.12 C 983.60,578.72 976.74,571.86 974.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1075.20,570.00 C 1064.22,580.98 1053.42,591.78 1050.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1024.80,570.00 C 1035.78,559.02 1046.58,548.22 1050.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,585.12 C 1043.60,578.72 1036.74,571.86 1034.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,554.88 C 1056.40,561.28 1063.26,568.14 1065.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1110.00,595.20 C 1099.02,584.22 1088.22,573.42 1084.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,544.80 C 1120.98,555.78 1131.78,566.58 1135.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1110.00,570.00 Q 1117.32,573.03 1123.20,570.00 Q 1117.32,566.97 1110.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,570.00 Q 1113.03,577.32 1119.33,579.33 Q 1117.32,573.03 1110.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,570.00 Q 1106.97,577.32 1110.00,583.20 Q 1113.03,577.32 1110.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,570.00 Q 1102.68,573.03 1100.67,579.33 Q 1106.97,577.32 1110.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,570.00 Q 1102.68,566.97 1096.80,570.00 Q 1102.68,573.03 1110.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,570.00 Q 1106.97,562.68 1100.67,560.67 Q 1102.68,566.97 1110.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,570.00 Q 1113.03,562.68 1110.00,556.80 Q 1106.97,562.68 1110.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,570.00 Q 1117.32,566.97 1119.33,560.67 Q 1113.03,562.68 1110.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,570.00 Q 1110.93,573.48 1115.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,570.00 Q 1106.52,570.93 1104.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,570.00 Q 1109.07,566.52 1104.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,570.00 Q 1113.48,569.07 1115.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1110.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1094.88,570.00 C 1101.28,563.60 1108.14,556.74 1110.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1125.12,570.00 C 1118.72,576.40 1111.86,583.26 1110.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1170.00,544.80 C 1180.98,555.78 1191.78,566.58 1195.20,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,595.20 C 1159.02,584.22 1148.22,573.42 1144.80,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1170.00,570.00 Q 1177.32,573.03 1183.20,570.00 Q 1177.32,566.97 1170.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,570.00 Q 1173.03,577.32 1179.33,579.33 Q 1177.32,573.03 1170.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,570.00 Q 1166.97,577.32 1170.00,583.20 Q 1173.03,577.32 1170.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,570.00 Q 1162.68,573.03 1160.67,579.33 Q 1166.97,577.32 1170.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,570.00 Q 1162.68,566.97 1156.80,570.00 Q 1162.68,573.03 1170.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,570.00 Q 1166.97,562.68 1160.67,560.67 Q 1162.68,566.97 1170.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,570.00 Q 1173.03,562.68 1170.00,556.80 Q 1166.97,562.68 1170.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,570.00 Q 1177.32,566.97 1179.33,560.67 Q 1173.03,562.68 1170.00,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,570.00 Q 1170.93,573.48 1175.09,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,570.00 Q 1166.52,570.93 1164.91,575.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,570.00 Q 1169.07,566.52 1164.91,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,570.00 Q 1173.48,569.07 1175.09,564.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1170.0" cy="570.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1185.12,570.00 C 1178.72,576.40 1171.86,583.26 1170.00,585.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1154.88,570.00 C 1161.28,563.60 1168.14,556.74 1170.00,554.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1204.80,570.00 C 1215.78,559.02 1226.58,548.22 1230.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1255.20,570.00 C 1244.22,580.98 1233.42,591.78 1230.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1230.00,554.88 C 1236.40,561.28 1243.26,568.14 1245.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,585.12 C 1223.60,578.72 1216.74,571.86 1214.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1315.20,570.00 C 1304.22,580.98 1293.42,591.78 1290.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1264.80,570.00 C 1275.78,559.02 1286.58,548.22 1290.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1290.00,585.12 C 1283.60,578.72 1276.74,571.86 1274.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,554.88 C 1296.40,561.28 1303.26,568.14 1305.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1324.80,570.00 C 1335.78,559.02 1346.58,548.22 1350.00,544.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1375.20,570.00 C 1364.22,580.98 1353.42,591.78 1350.00,595.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,554.88 C 1356.40,561.28 1363.26,568.14 1365.12,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,585.12 C 1343.60,578.72 1336.74,571.86 1334.88,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,604.80 C 160.98,615.78 171.78,626.58 175.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,655.20 C 139.02,644.22 128.22,633.42 124.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,630.00 Q 157.32,633.03 163.20,630.00 Q 157.32,626.97 150.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,630.00 Q 153.03,637.32 159.33,639.33 Q 157.32,633.03 150.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,630.00 Q 146.97,637.32 150.00,643.20 Q 153.03,637.32 150.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,630.00 Q 142.68,633.03 140.67,639.33 Q 146.97,637.32 150.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,630.00 Q 142.68,626.97 136.80,630.00 Q 142.68,633.03 150.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,630.00 Q 146.97,622.68 140.67,620.67 Q 142.68,626.97 150.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,630.00 Q 153.03,622.68 150.00,616.80 Q 146.97,622.68 150.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,630.00 Q 157.32,626.97 159.33,620.67 Q 153.03,622.68 150.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,630.00 Q 150.93,633.48 155.09,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,630.00 Q 146.52,630.93 144.91,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,630.00 Q 149.07,626.52 144.91,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,630.00 Q 153.48,629.07 155.09,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="630.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 165.12,630.00 C 158.72,636.40 151.86,643.26 150.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 134.88,630.00 C 141.28,623.60 148.14,616.74 150.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 235.20,630.00 C 224.22,640.98 213.42,651.78 210.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 184.80,630.00 C 195.78,619.02 206.58,608.22 210.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 210.00,630.00 Q 217.32,633.03 223.20,630.00 Q 217.32,626.97 210.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,630.00 Q 213.03,637.32 219.33,639.33 Q 217.32,633.03 210.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,630.00 Q 206.97,637.32 210.00,643.20 Q 213.03,637.32 210.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,630.00 Q 202.68,633.03 200.67,639.33 Q 206.97,637.32 210.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,630.00 Q 202.68,626.97 196.80,630.00 Q 202.68,633.03 210.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,630.00 Q 206.97,622.68 200.67,620.67 Q 202.68,626.97 210.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,630.00 Q 213.03,622.68 210.00,616.80 Q 206.97,622.68 210.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,630.00 Q 217.32,626.97 219.33,620.67 Q 213.03,622.68 210.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,630.00 Q 210.93,633.48 215.09,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,630.00 Q 206.52,630.93 204.91,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,630.00 Q 209.07,626.52 204.91,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,630.00 Q 213.48,629.07 215.09,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="210.0" cy="630.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 210.00,645.12 C 203.60,638.72 196.74,631.86 194.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,614.88 C 216.40,621.28 223.26,628.14 225.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,655.20 C 259.02,644.22 248.22,633.42 244.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,604.80 C 280.98,615.78 291.78,626.58 295.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 254.88,630.00 C 261.28,623.60 268.14,616.74 270.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 285.12,630.00 C 278.72,636.40 271.86,643.26 270.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 330.00,655.20 C 319.02,644.22 308.22,633.42 304.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,604.80 C 340.98,615.78 351.78,626.58 355.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 314.88,630.00 C 321.28,623.60 328.14,616.74 330.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 345.12,630.00 C 338.72,636.40 331.86,643.26 330.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 390.00,604.80 C 400.98,615.78 411.78,626.58 415.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,655.20 C 379.02,644.22 368.22,633.42 364.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 405.12,630.00 C 398.72,636.40 391.86,643.26 390.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 374.88,630.00 C 381.28,623.60 388.14,616.74 390.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 475.20,630.00 C 464.22,640.98 453.42,651.78 450.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 424.80,630.00 C 435.78,619.02 446.58,608.22 450.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 450.00,630.00 Q 457.32,633.03 463.20,630.00 Q 457.32,626.97 450.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,630.00 Q 453.03,637.32 459.33,639.33 Q 457.32,633.03 450.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,630.00 Q 446.97,637.32 450.00,643.20 Q 453.03,637.32 450.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,630.00 Q 442.68,633.03 440.67,639.33 Q 446.97,637.32 450.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,630.00 Q 442.68,626.97 436.80,630.00 Q 442.68,633.03 450.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,630.00 Q 446.97,622.68 440.67,620.67 Q 442.68,626.97 450.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,630.00 Q 453.03,622.68 450.00,616.80 Q 446.97,622.68 450.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,630.00 Q 457.32,626.97 459.33,620.67 Q 453.03,622.68 450.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,630.00 Q 450.93,633.48 455.09,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,630.00 Q 446.52,630.93 444.91,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,630.00 Q 449.07,626.52 444.91,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,630.00 Q 453.48,629.07 455.09,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="450.0" cy="630.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 450.00,645.12 C 443.60,638.72 436.74,631.86 434.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,614.88 C 456.40,621.28 463.26,628.14 465.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 535.20,630.00 C 524.22,640.98 513.42,651.78 510.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 484.80,630.00 C 495.78,619.02 506.58,608.22 510.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,630.00 Q 517.32,633.03 523.20,630.00 Q 517.32,626.97 510.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,630.00 Q 513.03,637.32 519.33,639.33 Q 517.32,633.03 510.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,630.00 Q 506.97,637.32 510.00,643.20 Q 513.03,637.32 510.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,630.00 Q 502.68,633.03 500.67,639.33 Q 506.97,637.32 510.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,630.00 Q 502.68,626.97 496.80,630.00 Q 502.68,633.03 510.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,630.00 Q 506.97,622.68 500.67,620.67 Q 502.68,626.97 510.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,630.00 Q 513.03,622.68 510.00,616.80 Q 506.97,622.68 510.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,630.00 Q 517.32,626.97 519.33,620.67 Q 513.03,622.68 510.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,630.00 Q 510.93,633.48 515.09,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,630.00 Q 506.52,630.93 504.91,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,630.00 Q 509.07,626.52 504.91,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,630.00 Q 513.48,629.07 515.09,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="630.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 510.00,645.12 C 503.60,638.72 496.74,631.86 494.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,614.88 C 516.40,621.28 523.26,628.14 525.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 570.00,655.20 C 559.02,644.22 548.22,633.42 544.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,604.80 C 580.98,615.78 591.78,626.58 595.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 554.88,630.00 C 561.28,623.60 568.14,616.74 570.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 585.12,630.00 C 578.72,636.40 571.86,643.26 570.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 630.00,604.80 C 640.98,615.78 651.78,626.58 655.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,655.20 C 619.02,644.22 608.22,633.42 604.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 630.00,630.00 Q 637.32,633.03 643.20,630.00 Q 637.32,626.97 630.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,630.00 Q 633.03,637.32 639.33,639.33 Q 637.32,633.03 630.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,630.00 Q 626.97,637.32 630.00,643.20 Q 633.03,637.32 630.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,630.00 Q 622.68,633.03 620.67,639.33 Q 626.97,637.32 630.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,630.00 Q 622.68,626.97 616.80,630.00 Q 622.68,633.03 630.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,630.00 Q 626.97,622.68 620.67,620.67 Q 622.68,626.97 630.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,630.00 Q 633.03,622.68 630.00,616.80 Q 626.97,622.68 630.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,630.00 Q 637.32,626.97 639.33,620.67 Q 633.03,622.68 630.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,630.00 Q 630.93,633.48 635.09,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,630.00 Q 626.52,630.93 624.91,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,630.00 Q 629.07,626.52 624.91,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,630.00 Q 633.48,629.07 635.09,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="630.0" cy="630.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 645.12,630.00 C 638.72,636.40 631.86,643.26 630.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 614.88,630.00 C 621.28,623.60 628.14,616.74 630.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 715.20,630.00 C 704.22,640.98 693.42,651.78 690.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 664.80,630.00 C 675.78,619.02 686.58,608.22 690.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 690.00,630.00 Q 697.32,633.03 703.20,630.00 Q 697.32,626.97 690.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,630.00 Q 693.03,637.32 699.33,639.33 Q 697.32,633.03 690.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,630.00 Q 686.97,637.32 690.00,643.20 Q 693.03,637.32 690.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,630.00 Q 682.68,633.03 680.67,639.33 Q 686.97,637.32 690.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,630.00 Q 682.68,626.97 676.80,630.00 Q 682.68,633.03 690.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,630.00 Q 686.97,622.68 680.67,620.67 Q 682.68,626.97 690.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,630.00 Q 693.03,622.68 690.00,616.80 Q 686.97,622.68 690.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,630.00 Q 697.32,626.97 699.33,620.67 Q 693.03,622.68 690.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,630.00 Q 690.93,633.48 695.09,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,630.00 Q 686.52,630.93 684.91,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,630.00 Q 689.07,626.52 684.91,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,630.00 Q 693.48,629.07 695.09,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="690.0" cy="630.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 690.00,645.12 C 683.60,638.72 676.74,631.86 674.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,614.88 C 696.40,621.28 703.26,628.14 705.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 775.20,630.00 C 764.22,640.98 753.42,651.78 750.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 724.80,630.00 C 735.78,619.02 746.58,608.22 750.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,645.12 C 743.60,638.72 736.74,631.86 734.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,614.88 C 756.40,621.28 763.26,628.14 765.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 810.00,655.20 C 799.02,644.22 788.22,633.42 784.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,604.80 C 820.98,615.78 831.78,626.58 835.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 794.88,630.00 C 801.28,623.60 808.14,616.74 810.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 825.12,630.00 C 818.72,636.40 811.86,643.26 810.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 895.20,630.00 C 884.22,640.98 873.42,651.78 870.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 844.80,630.00 C 855.78,619.02 866.58,608.22 870.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,630.00 Q 877.32,633.03 883.20,630.00 Q 877.32,626.97 870.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,630.00 Q 873.03,637.32 879.33,639.33 Q 877.32,633.03 870.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,630.00 Q 866.97,637.32 870.00,643.20 Q 873.03,637.32 870.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,630.00 Q 862.68,633.03 860.67,639.33 Q 866.97,637.32 870.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,630.00 Q 862.68,626.97 856.80,630.00 Q 862.68,633.03 870.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,630.00 Q 866.97,622.68 860.67,620.67 Q 862.68,626.97 870.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,630.00 Q 873.03,622.68 870.00,616.80 Q 866.97,622.68 870.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,630.00 Q 877.32,626.97 879.33,620.67 Q 873.03,622.68 870.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,630.00 Q 870.93,633.48 875.09,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,630.00 Q 866.52,630.93 864.91,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,630.00 Q 869.07,626.52 864.91,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,630.00 Q 873.48,629.07 875.09,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="630.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 870.00,645.12 C 863.60,638.72 856.74,631.86 854.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,614.88 C 876.40,621.28 883.26,628.14 885.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 955.20,630.00 C 944.22,640.98 933.42,651.78 930.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 904.80,630.00 C 915.78,619.02 926.58,608.22 930.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,630.00 Q 937.32,633.03 943.20,630.00 Q 937.32,626.97 930.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,630.00 Q 933.03,637.32 939.33,639.33 Q 937.32,633.03 930.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,630.00 Q 926.97,637.32 930.00,643.20 Q 933.03,637.32 930.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,630.00 Q 922.68,633.03 920.67,639.33 Q 926.97,637.32 930.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,630.00 Q 922.68,626.97 916.80,630.00 Q 922.68,633.03 930.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,630.00 Q 926.97,622.68 920.67,620.67 Q 922.68,626.97 930.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,630.00 Q 933.03,622.68 930.00,616.80 Q 926.97,622.68 930.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,630.00 Q 937.32,626.97 939.33,620.67 Q 933.03,622.68 930.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,630.00 Q 930.93,633.48 935.09,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,630.00 Q 926.52,630.93 924.91,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,630.00 Q 929.07,626.52 924.91,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,630.00 Q 933.48,629.07 935.09,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="630.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 930.00,645.12 C 923.60,638.72 916.74,631.86 914.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,614.88 C 936.40,621.28 943.26,628.14 945.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,655.20 C 979.02,644.22 968.22,633.42 964.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,604.80 C 1000.98,615.78 1011.78,626.58 1015.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 974.88,630.00 C 981.28,623.60 988.14,616.74 990.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1005.12,630.00 C 998.72,636.40 991.86,643.26 990.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1050.00,655.20 C 1039.02,644.22 1028.22,633.42 1024.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,604.80 C 1060.98,615.78 1071.78,626.58 1075.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1034.88,630.00 C 1041.28,623.60 1048.14,616.74 1050.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1065.12,630.00 C 1058.72,636.40 1051.86,643.26 1050.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1084.80,630.00 C 1095.78,619.02 1106.58,608.22 1110.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1135.20,630.00 C 1124.22,640.98 1113.42,651.78 1110.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1110.00,630.00 Q 1117.32,633.03 1123.20,630.00 Q 1117.32,626.97 1110.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,630.00 Q 1113.03,637.32 1119.33,639.33 Q 1117.32,633.03 1110.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,630.00 Q 1106.97,637.32 1110.00,643.20 Q 1113.03,637.32 1110.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,630.00 Q 1102.68,633.03 1100.67,639.33 Q 1106.97,637.32 1110.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,630.00 Q 1102.68,626.97 1096.80,630.00 Q 1102.68,633.03 1110.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,630.00 Q 1106.97,622.68 1100.67,620.67 Q 1102.68,626.97 1110.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,630.00 Q 1113.03,622.68 1110.00,616.80 Q 1106.97,622.68 1110.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,630.00 Q 1117.32,626.97 1119.33,620.67 Q 1113.03,622.68 1110.00,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,630.00 Q 1110.93,633.48 1115.09,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,630.00 Q 1106.52,630.93 1104.91,635.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,630.00 Q 1109.07,626.52 1104.91,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,630.00 Q 1113.48,629.07 1115.09,624.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1110.0" cy="630.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1110.00,614.88 C 1116.40,621.28 1123.26,628.14 1125.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,645.12 C 1103.60,638.72 1096.74,631.86 1094.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1144.80,630.00 C 1155.78,619.02 1166.58,608.22 1170.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1195.20,630.00 C 1184.22,640.98 1173.42,651.78 1170.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1170.00,614.88 C 1176.40,621.28 1183.26,628.14 1185.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,645.12 C 1163.60,638.72 1156.74,631.86 1154.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1204.80,630.00 C 1215.78,619.02 1226.58,608.22 1230.00,604.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1255.20,630.00 C 1244.22,640.98 1233.42,651.78 1230.00,655.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1230.00,614.88 C 1236.40,621.28 1243.26,628.14 1245.12,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,645.12 C 1223.60,638.72 1216.74,631.86 1214.88,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1290.00,655.20 C 1279.02,644.22 1268.22,633.42 1264.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,604.80 C 1300.98,615.78 1311.78,626.58 1315.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1274.88,630.00 C 1281.28,623.60 1288.14,616.74 1290.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1305.12,630.00 C 1298.72,636.40 1291.86,643.26 1290.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1350.00,604.80 C 1360.98,615.78 1371.78,626.58 1375.20,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,655.20 C 1339.02,644.22 1328.22,633.42 1324.80,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1365.12,630.00 C 1358.72,636.40 1351.86,643.26 1350.00,645.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1334.88,630.00 C 1341.28,623.60 1348.14,616.74 1350.00,614.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 175.20,690.00 C 164.22,700.98 153.42,711.78 150.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 124.80,690.00 C 135.78,679.02 146.58,668.22 150.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,690.00 Q 157.32,693.03 163.20,690.00 Q 157.32,686.97 150.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,690.00 Q 153.03,697.32 159.33,699.33 Q 157.32,693.03 150.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,690.00 Q 146.97,697.32 150.00,703.20 Q 153.03,697.32 150.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,690.00 Q 142.68,693.03 140.67,699.33 Q 146.97,697.32 150.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,690.00 Q 142.68,686.97 136.80,690.00 Q 142.68,693.03 150.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,690.00 Q 146.97,682.68 140.67,680.67 Q 142.68,686.97 150.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,690.00 Q 153.03,682.68 150.00,676.80 Q 146.97,682.68 150.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,690.00 Q 157.32,686.97 159.33,680.67 Q 153.03,682.68 150.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,690.00 Q 150.93,693.48 155.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,690.00 Q 146.52,690.93 144.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,690.00 Q 149.07,686.52 144.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,690.00 Q 153.48,689.07 155.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 150.00,705.12 C 143.60,698.72 136.74,691.86 134.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,674.88 C 156.40,681.28 163.26,688.14 165.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 235.20,690.00 C 224.22,700.98 213.42,711.78 210.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 184.80,690.00 C 195.78,679.02 206.58,668.22 210.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 210.00,690.00 Q 217.32,693.03 223.20,690.00 Q 217.32,686.97 210.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,690.00 Q 213.03,697.32 219.33,699.33 Q 217.32,693.03 210.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,690.00 Q 206.97,697.32 210.00,703.20 Q 213.03,697.32 210.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,690.00 Q 202.68,693.03 200.67,699.33 Q 206.97,697.32 210.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,690.00 Q 202.68,686.97 196.80,690.00 Q 202.68,693.03 210.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,690.00 Q 206.97,682.68 200.67,680.67 Q 202.68,686.97 210.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,690.00 Q 213.03,682.68 210.00,676.80 Q 206.97,682.68 210.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,690.00 Q 217.32,686.97 219.33,680.67 Q 213.03,682.68 210.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,690.00 Q 210.93,693.48 215.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,690.00 Q 206.52,690.93 204.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,690.00 Q 209.07,686.52 204.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,690.00 Q 213.48,689.07 215.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="210.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 210.00,705.12 C 203.60,698.72 196.74,691.86 194.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,674.88 C 216.40,681.28 223.26,688.14 225.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,664.80 C 280.98,675.78 291.78,686.58 295.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,715.20 C 259.02,704.22 248.22,693.42 244.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 270.00,690.00 Q 277.32,693.03 283.20,690.00 Q 277.32,686.97 270.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,690.00 Q 273.03,697.32 279.33,699.33 Q 277.32,693.03 270.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,690.00 Q 266.97,697.32 270.00,703.20 Q 273.03,697.32 270.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,690.00 Q 262.68,693.03 260.67,699.33 Q 266.97,697.32 270.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,690.00 Q 262.68,686.97 256.80,690.00 Q 262.68,693.03 270.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,690.00 Q 266.97,682.68 260.67,680.67 Q 262.68,686.97 270.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,690.00 Q 273.03,682.68 270.00,676.80 Q 266.97,682.68 270.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,690.00 Q 277.32,686.97 279.33,680.67 Q 273.03,682.68 270.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,690.00 Q 270.93,693.48 275.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,690.00 Q 266.52,690.93 264.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,690.00 Q 269.07,686.52 264.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,690.00 Q 273.48,689.07 275.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="270.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 285.12,690.00 C 278.72,696.40 271.86,703.26 270.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 254.88,690.00 C 261.28,683.60 268.14,676.74 270.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 330.00,664.80 C 340.98,675.78 351.78,686.58 355.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,715.20 C 319.02,704.22 308.22,693.42 304.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 330.00,690.00 Q 337.32,693.03 343.20,690.00 Q 337.32,686.97 330.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,690.00 Q 333.03,697.32 339.33,699.33 Q 337.32,693.03 330.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,690.00 Q 326.97,697.32 330.00,703.20 Q 333.03,697.32 330.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,690.00 Q 322.68,693.03 320.67,699.33 Q 326.97,697.32 330.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,690.00 Q 322.68,686.97 316.80,690.00 Q 322.68,693.03 330.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,690.00 Q 326.97,682.68 320.67,680.67 Q 322.68,686.97 330.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,690.00 Q 333.03,682.68 330.00,676.80 Q 326.97,682.68 330.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,690.00 Q 337.32,686.97 339.33,680.67 Q 333.03,682.68 330.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,690.00 Q 330.93,693.48 335.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,690.00 Q 326.52,690.93 324.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,690.00 Q 329.07,686.52 324.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,690.00 Q 333.48,689.07 335.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="330.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 345.12,690.00 C 338.72,696.40 331.86,703.26 330.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 314.88,690.00 C 321.28,683.60 328.14,676.74 330.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 415.20,690.00 C 404.22,700.98 393.42,711.78 390.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 364.80,690.00 C 375.78,679.02 386.58,668.22 390.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 390.00,690.00 Q 397.32,693.03 403.20,690.00 Q 397.32,686.97 390.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,690.00 Q 393.03,697.32 399.33,699.33 Q 397.32,693.03 390.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,690.00 Q 386.97,697.32 390.00,703.20 Q 393.03,697.32 390.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,690.00 Q 382.68,693.03 380.67,699.33 Q 386.97,697.32 390.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,690.00 Q 382.68,686.97 376.80,690.00 Q 382.68,693.03 390.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,690.00 Q 386.97,682.68 380.67,680.67 Q 382.68,686.97 390.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,690.00 Q 393.03,682.68 390.00,676.80 Q 386.97,682.68 390.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,690.00 Q 397.32,686.97 399.33,680.67 Q 393.03,682.68 390.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,690.00 Q 390.93,693.48 395.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,690.00 Q 386.52,690.93 384.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,690.00 Q 389.07,686.52 384.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,690.00 Q 393.48,689.07 395.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="390.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 390.00,705.12 C 383.60,698.72 376.74,691.86 374.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,674.88 C 396.40,681.28 403.26,688.14 405.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 475.20,690.00 C 464.22,700.98 453.42,711.78 450.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 424.80,690.00 C 435.78,679.02 446.58,668.22 450.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 450.00,705.12 C 443.60,698.72 436.74,691.86 434.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,674.88 C 456.40,681.28 463.26,688.14 465.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,715.20 C 499.02,704.22 488.22,693.42 484.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,664.80 C 520.98,675.78 531.78,686.58 535.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 494.88,690.00 C 501.28,683.60 508.14,676.74 510.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 525.12,690.00 C 518.72,696.40 511.86,703.26 510.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 570.00,664.80 C 580.98,675.78 591.78,686.58 595.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,715.20 C 559.02,704.22 548.22,693.42 544.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 585.12,690.00 C 578.72,696.40 571.86,703.26 570.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 554.88,690.00 C 561.28,683.60 568.14,676.74 570.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 655.20,690.00 C 644.22,700.98 633.42,711.78 630.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 604.80,690.00 C 615.78,679.02 626.58,668.22 630.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,705.12 C 623.60,698.72 616.74,691.86 614.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,674.88 C 636.40,681.28 643.26,688.14 645.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 715.20,690.00 C 704.22,700.98 693.42,711.78 690.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 664.80,690.00 C 675.78,679.02 686.58,668.22 690.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 690.00,705.12 C 683.60,698.72 676.74,691.86 674.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,674.88 C 696.40,681.28 703.26,688.14 705.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 724.80,690.00 C 735.78,679.02 746.58,668.22 750.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 775.20,690.00 C 764.22,700.98 753.42,711.78 750.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,674.88 C 756.40,681.28 763.26,688.14 765.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,705.12 C 743.60,698.72 736.74,691.86 734.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 810.00,664.80 C 820.98,675.78 831.78,686.58 835.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,715.20 C 799.02,704.22 788.22,693.42 784.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 810.00,690.00 Q 817.32,693.03 823.20,690.00 Q 817.32,686.97 810.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,690.00 Q 813.03,697.32 819.33,699.33 Q 817.32,693.03 810.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,690.00 Q 806.97,697.32 810.00,703.20 Q 813.03,697.32 810.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,690.00 Q 802.68,693.03 800.67,699.33 Q 806.97,697.32 810.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,690.00 Q 802.68,686.97 796.80,690.00 Q 802.68,693.03 810.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,690.00 Q 806.97,682.68 800.67,680.67 Q 802.68,686.97 810.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,690.00 Q 813.03,682.68 810.00,676.80 Q 806.97,682.68 810.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,690.00 Q 817.32,686.97 819.33,680.67 Q 813.03,682.68 810.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,690.00 Q 810.93,693.48 815.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,690.00 Q 806.52,690.93 804.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,690.00 Q 809.07,686.52 804.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,690.00 Q 813.48,689.07 815.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="810.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 825.12,690.00 C 818.72,696.40 811.86,703.26 810.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 794.88,690.00 C 801.28,683.60 808.14,676.74 810.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 895.20,690.00 C 884.22,700.98 873.42,711.78 870.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 844.80,690.00 C 855.78,679.02 866.58,668.22 870.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,690.00 Q 877.32,693.03 883.20,690.00 Q 877.32,686.97 870.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,690.00 Q 873.03,697.32 879.33,699.33 Q 877.32,693.03 870.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,690.00 Q 866.97,697.32 870.00,703.20 Q 873.03,697.32 870.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,690.00 Q 862.68,693.03 860.67,699.33 Q 866.97,697.32 870.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,690.00 Q 862.68,686.97 856.80,690.00 Q 862.68,693.03 870.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,690.00 Q 866.97,682.68 860.67,680.67 Q 862.68,686.97 870.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,690.00 Q 873.03,682.68 870.00,676.80 Q 866.97,682.68 870.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,690.00 Q 877.32,686.97 879.33,680.67 Q 873.03,682.68 870.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,690.00 Q 870.93,693.48 875.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,690.00 Q 866.52,690.93 864.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,690.00 Q 869.07,686.52 864.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,690.00 Q 873.48,689.07 875.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 870.00,705.12 C 863.60,698.72 856.74,691.86 854.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,674.88 C 876.40,681.28 883.26,688.14 885.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 930.00,715.20 C 919.02,704.22 908.22,693.42 904.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,664.80 C 940.98,675.78 951.78,686.58 955.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 914.88,690.00 C 921.28,683.60 928.14,676.74 930.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 945.12,690.00 C 938.72,696.40 931.86,703.26 930.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,715.20 C 979.02,704.22 968.22,693.42 964.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,664.80 C 1000.98,675.78 1011.78,686.58 1015.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 974.88,690.00 C 981.28,683.60 988.14,676.74 990.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1005.12,690.00 C 998.72,696.40 991.86,703.26 990.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1075.20,690.00 C 1064.22,700.98 1053.42,711.78 1050.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1024.80,690.00 C 1035.78,679.02 1046.58,668.22 1050.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1050.00,690.00 Q 1057.32,693.03 1063.20,690.00 Q 1057.32,686.97 1050.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,690.00 Q 1053.03,697.32 1059.33,699.33 Q 1057.32,693.03 1050.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,690.00 Q 1046.97,697.32 1050.00,703.20 Q 1053.03,697.32 1050.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,690.00 Q 1042.68,693.03 1040.67,699.33 Q 1046.97,697.32 1050.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,690.00 Q 1042.68,686.97 1036.80,690.00 Q 1042.68,693.03 1050.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,690.00 Q 1046.97,682.68 1040.67,680.67 Q 1042.68,686.97 1050.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,690.00 Q 1053.03,682.68 1050.00,676.80 Q 1046.97,682.68 1050.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,690.00 Q 1057.32,686.97 1059.33,680.67 Q 1053.03,682.68 1050.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,690.00 Q 1050.93,693.48 1055.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,690.00 Q 1046.52,690.93 1044.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,690.00 Q 1049.07,686.52 1044.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,690.00 Q 1053.48,689.07 1055.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1050.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1050.00,705.12 C 1043.60,698.72 1036.74,691.86 1034.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,674.88 C 1056.40,681.28 1063.26,688.14 1065.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1135.20,690.00 C 1124.22,700.98 1113.42,711.78 1110.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1084.80,690.00 C 1095.78,679.02 1106.58,668.22 1110.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1110.00,690.00 Q 1117.32,693.03 1123.20,690.00 Q 1117.32,686.97 1110.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,690.00 Q 1113.03,697.32 1119.33,699.33 Q 1117.32,693.03 1110.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,690.00 Q 1106.97,697.32 1110.00,703.20 Q 1113.03,697.32 1110.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,690.00 Q 1102.68,693.03 1100.67,699.33 Q 1106.97,697.32 1110.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,690.00 Q 1102.68,686.97 1096.80,690.00 Q 1102.68,693.03 1110.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,690.00 Q 1106.97,682.68 1100.67,680.67 Q 1102.68,686.97 1110.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,690.00 Q 1113.03,682.68 1110.00,676.80 Q 1106.97,682.68 1110.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,690.00 Q 1117.32,686.97 1119.33,680.67 Q 1113.03,682.68 1110.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,690.00 Q 1110.93,693.48 1115.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,690.00 Q 1106.52,690.93 1104.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,690.00 Q 1109.07,686.52 1104.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,690.00 Q 1113.48,689.07 1115.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1110.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1110.00,705.12 C 1103.60,698.72 1096.74,691.86 1094.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,674.88 C 1116.40,681.28 1123.26,688.14 1125.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1170.00,715.20 C 1159.02,704.22 1148.22,693.42 1144.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,664.80 C 1180.98,675.78 1191.78,686.58 1195.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1154.88,690.00 C 1161.28,683.60 1168.14,676.74 1170.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1185.12,690.00 C 1178.72,696.40 1171.86,703.26 1170.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,715.20 C 1219.02,704.22 1208.22,693.42 1204.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,664.80 C 1240.98,675.78 1251.78,686.58 1255.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1230.00,690.00 Q 1237.32,693.03 1243.20,690.00 Q 1237.32,686.97 1230.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,690.00 Q 1233.03,697.32 1239.33,699.33 Q 1237.32,693.03 1230.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,690.00 Q 1226.97,697.32 1230.00,703.20 Q 1233.03,697.32 1230.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,690.00 Q 1222.68,693.03 1220.67,699.33 Q 1226.97,697.32 1230.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,690.00 Q 1222.68,686.97 1216.80,690.00 Q 1222.68,693.03 1230.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,690.00 Q 1226.97,682.68 1220.67,680.67 Q 1222.68,686.97 1230.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,690.00 Q 1233.03,682.68 1230.00,676.80 Q 1226.97,682.68 1230.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,690.00 Q 1237.32,686.97 1239.33,680.67 Q 1233.03,682.68 1230.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,690.00 Q 1230.93,693.48 1235.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,690.00 Q 1226.52,690.93 1224.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,690.00 Q 1229.07,686.52 1224.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,690.00 Q 1233.48,689.07 1235.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1230.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1214.88,690.00 C 1221.28,683.60 1228.14,676.74 1230.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1245.12,690.00 C 1238.72,696.40 1231.86,703.26 1230.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1290.00,664.80 C 1300.98,675.78 1311.78,686.58 1315.20,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,715.20 C 1279.02,704.22 1268.22,693.42 1264.80,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1290.00,690.00 Q 1297.32,693.03 1303.20,690.00 Q 1297.32,686.97 1290.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,690.00 Q 1293.03,697.32 1299.33,699.33 Q 1297.32,693.03 1290.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,690.00 Q 1286.97,697.32 1290.00,703.20 Q 1293.03,697.32 1290.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,690.00 Q 1282.68,693.03 1280.67,699.33 Q 1286.97,697.32 1290.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,690.00 Q 1282.68,686.97 1276.80,690.00 Q 1282.68,693.03 1290.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,690.00 Q 1286.97,682.68 1280.67,680.67 Q 1282.68,686.97 1290.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,690.00 Q 1293.03,682.68 1290.00,676.80 Q 1286.97,682.68 1290.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,690.00 Q 1297.32,686.97 1299.33,680.67 Q 1293.03,682.68 1290.00,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,690.00 Q 1290.93,693.48 1295.09,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,690.00 Q 1286.52,690.93 1284.91,695.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,690.00 Q 1289.07,686.52 1284.91,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,690.00 Q 1293.48,689.07 1295.09,684.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1290.0" cy="690.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1305.12,690.00 C 1298.72,696.40 1291.86,703.26 1290.00,705.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1274.88,690.00 C 1281.28,683.60 1288.14,676.74 1290.00,674.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1375.20,690.00 C 1364.22,700.98 1353.42,711.78 1350.00,715.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1324.80,690.00 C 1335.78,679.02 1346.58,668.22 1350.00,664.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,705.12 C 1343.60,698.72 1336.74,691.86 1334.88,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,674.88 C 1356.40,681.28 1363.26,688.14 1365.12,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,724.80 C 160.98,735.78 171.78,746.58 175.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,775.20 C 139.02,764.22 128.22,753.42 124.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 165.12,750.00 C 158.72,756.40 151.86,763.26 150.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 134.88,750.00 C 141.28,743.60 148.14,736.74 150.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 210.00,775.20 C 199.02,764.22 188.22,753.42 184.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,724.80 C 220.98,735.78 231.78,746.58 235.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 194.88,750.00 C 201.28,743.60 208.14,736.74 210.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 225.12,750.00 C 218.72,756.40 211.86,763.26 210.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,775.20 C 259.02,764.22 248.22,753.42 244.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,724.80 C 280.98,735.78 291.78,746.58 295.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 270.00,750.00 Q 277.32,753.03 283.20,750.00 Q 277.32,746.97 270.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,750.00 Q 273.03,757.32 279.33,759.33 Q 277.32,753.03 270.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,750.00 Q 266.97,757.32 270.00,763.20 Q 273.03,757.32 270.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,750.00 Q 262.68,753.03 260.67,759.33 Q 266.97,757.32 270.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,750.00 Q 262.68,746.97 256.80,750.00 Q 262.68,753.03 270.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,750.00 Q 266.97,742.68 260.67,740.67 Q 262.68,746.97 270.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,750.00 Q 273.03,742.68 270.00,736.80 Q 266.97,742.68 270.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,750.00 Q 277.32,746.97 279.33,740.67 Q 273.03,742.68 270.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,750.00 Q 270.93,753.48 275.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,750.00 Q 266.52,750.93 264.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,750.00 Q 269.07,746.52 264.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,750.00 Q 273.48,749.07 275.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="270.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 254.88,750.00 C 261.28,743.60 268.14,736.74 270.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 285.12,750.00 C 278.72,756.40 271.86,763.26 270.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 355.20,750.00 C 344.22,760.98 333.42,771.78 330.00,775.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 304.80,750.00 C 315.78,739.02 326.58,728.22 330.00,724.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 330.00,750.00 Q 337.32,753.03 343.20,750.00 Q 337.32,746.97 330.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,750.00 Q 333.03,757.32 339.33,759.33 Q 337.32,753.03 330.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,750.00 Q 326.97,757.32 330.00,763.20 Q 333.03,757.32 330.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,750.00 Q 322.68,753.03 320.67,759.33 Q 326.97,757.32 330.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,750.00 Q 322.68,746.97 316.80,750.00 Q 322.68,753.03 330.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,750.00 Q 326.97,742.68 320.67,740.67 Q 322.68,746.97 330.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,750.00 Q 333.03,742.68 330.00,736.80 Q 326.97,742.68 330.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,750.00 Q 337.32,746.97 339.33,740.67 Q 333.03,742.68 330.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,750.00 Q 330.93,753.48 335.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,750.00 Q 326.52,750.93 324.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,750.00 Q 329.07,746.52 324.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,750.00 Q 333.48,749.07 335.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="330.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 330.00,765.12 C 323.60,758.72 316.74,751.86 314.88,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,734.88 C 336.40,741.28 343.26,748.14 345.12,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 415.20,750.00 C 404.22,760.98 393.42,771.78 390.00,775.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 364.80,750.00 C 375.78,739.02 386.58,728.22 390.00,724.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 390.00,750.00 Q 397.32,753.03 403.20,750.00 Q 397.32,746.97 390.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,750.00 Q 393.03,757.32 399.33,759.33 Q 397.32,753.03 390.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,750.00 Q 386.97,757.32 390.00,763.20 Q 393.03,757.32 390.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,750.00 Q 382.68,753.03 380.67,759.33 Q 386.97,757.32 390.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,750.00 Q 382.68,746.97 376.80,750.00 Q 382.68,753.03 390.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,750.00 Q 386.97,742.68 380.67,740.67 Q 382.68,746.97 390.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,750.00 Q 393.03,742.68 390.00,736.80 Q 386.97,742.68 390.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,750.00 Q 397.32,746.97 399.33,740.67 Q 393.03,742.68 390.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,750.00 Q 390.93,753.48 395.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,750.00 Q 386.52,750.93 384.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,750.00 Q 389.07,746.52 384.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,750.00 Q 393.48,749.07 395.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="390.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 390.00,765.12 C 383.60,758.72 376.74,751.86 374.88,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,734.88 C 396.40,741.28 403.26,748.14 405.12,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 450.00,724.80 C 460.98,735.78 471.78,746.58 475.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,775.20 C 439.02,764.22 428.22,753.42 424.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 465.12,750.00 C 458.72,756.40 451.86,763.26 450.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 434.88,750.00 C 441.28,743.60 448.14,736.74 450.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,724.80 C 520.98,735.78 531.78,746.58 535.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,775.20 C 499.02,764.22 488.22,753.42 484.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,750.00 Q 517.32,753.03 523.20,750.00 Q 517.32,746.97 510.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,750.00 Q 513.03,757.32 519.33,759.33 Q 517.32,753.03 510.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,750.00 Q 506.97,757.32 510.00,763.20 Q 513.03,757.32 510.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,750.00 Q 502.68,753.03 500.67,759.33 Q 506.97,757.32 510.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,750.00 Q 502.68,746.97 496.80,750.00 Q 502.68,753.03 510.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,750.00 Q 506.97,742.68 500.67,740.67 Q 502.68,746.97 510.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,750.00 Q 513.03,742.68 510.00,736.80 Q 506.97,742.68 510.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,750.00 Q 517.32,746.97 519.33,740.67 Q 513.03,742.68 510.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,750.00 Q 510.93,753.48 515.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,750.00 Q 506.52,750.93 504.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,750.00 Q 509.07,746.52 504.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,750.00 Q 513.48,749.07 515.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 525.12,750.00 C 518.72,756.40 511.86,763.26 510.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 494.88,750.00 C 501.28,743.60 508.14,736.74 510.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,750.00 C 555.78,739.02 566.58,728.22 570.00,724.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,750.00 C 584.22,760.98 573.42,771.78 570.00,775.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 570.00,750.00 Q 577.32,753.03 583.20,750.00 Q 577.32,746.97 570.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,750.00 Q 573.03,757.32 579.33,759.33 Q 577.32,753.03 570.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,750.00 Q 566.97,757.32 570.00,763.20 Q 573.03,757.32 570.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,750.00 Q 562.68,753.03 560.67,759.33 Q 566.97,757.32 570.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,750.00 Q 562.68,746.97 556.80,750.00 Q 562.68,753.03 570.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,750.00 Q 566.97,742.68 560.67,740.67 Q 562.68,746.97 570.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,750.00 Q 573.03,742.68 570.00,736.80 Q 566.97,742.68 570.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,750.00 Q 577.32,746.97 579.33,740.67 Q 573.03,742.68 570.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,750.00 Q 570.93,753.48 575.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,750.00 Q 566.52,750.93 564.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,750.00 Q 569.07,746.52 564.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,750.00 Q 573.48,749.07 575.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="570.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 570.00,734.88 C 576.40,741.28 583.26,748.14 585.12,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,765.12 C 563.60,758.72 556.74,751.86 554.88,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 630.00,724.80 C 640.98,735.78 651.78,746.58 655.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,775.20 C 619.02,764.22 608.22,753.42 604.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 645.12,750.00 C 638.72,756.40 631.86,763.26 630.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 614.88,750.00 C 621.28,743.60 628.14,736.74 630.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 690.00,775.20 C 679.02,764.22 668.22,753.42 664.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,724.80 C 700.98,735.78 711.78,746.58 715.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 674.88,750.00 C 681.28,743.60 688.14,736.74 690.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 705.12,750.00 C 698.72,756.40 691.86,763.26 690.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 775.20,750.00 C 764.22,760.98 753.42,771.78 750.00,775.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 724.80,750.00 C 735.78,739.02 746.58,728.22 750.00,724.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 750.00,750.00 Q 757.32,753.03 763.20,750.00 Q 757.32,746.97 750.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,750.00 Q 753.03,757.32 759.33,759.33 Q 757.32,753.03 750.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,750.00 Q 746.97,757.32 750.00,763.20 Q 753.03,757.32 750.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,750.00 Q 742.68,753.03 740.67,759.33 Q 746.97,757.32 750.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,750.00 Q 742.68,746.97 736.80,750.00 Q 742.68,753.03 750.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,750.00 Q 746.97,742.68 740.67,740.67 Q 742.68,746.97 750.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,750.00 Q 753.03,742.68 750.00,736.80 Q 746.97,742.68 750.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,750.00 Q 757.32,746.97 759.33,740.67 Q 753.03,742.68 750.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,750.00 Q 750.93,753.48 755.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,750.00 Q 746.52,750.93 744.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,750.00 Q 749.07,746.52 744.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,750.00 Q 753.48,749.07 755.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="750.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 750.00,765.12 C 743.60,758.72 736.74,751.86 734.88,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,734.88 C 756.40,741.28 763.26,748.14 765.12,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 835.20,750.00 C 824.22,760.98 813.42,771.78 810.00,775.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 784.80,750.00 C 795.78,739.02 806.58,728.22 810.00,724.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 810.00,750.00 Q 817.32,753.03 823.20,750.00 Q 817.32,746.97 810.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,750.00 Q 813.03,757.32 819.33,759.33 Q 817.32,753.03 810.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,750.00 Q 806.97,757.32 810.00,763.20 Q 813.03,757.32 810.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,750.00 Q 802.68,753.03 800.67,759.33 Q 806.97,757.32 810.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,750.00 Q 802.68,746.97 796.80,750.00 Q 802.68,753.03 810.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,750.00 Q 806.97,742.68 800.67,740.67 Q 802.68,746.97 810.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,750.00 Q 813.03,742.68 810.00,736.80 Q 806.97,742.68 810.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,750.00 Q 817.32,746.97 819.33,740.67 Q 813.03,742.68 810.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,750.00 Q 810.93,753.48 815.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,750.00 Q 806.52,750.93 804.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,750.00 Q 809.07,746.52 804.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,750.00 Q 813.48,749.07 815.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="810.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 810.00,765.12 C 803.60,758.72 796.74,751.86 794.88,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,734.88 C 816.40,741.28 823.26,748.14 825.12,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 870.00,775.20 C 859.02,764.22 848.22,753.42 844.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,724.80 C 880.98,735.78 891.78,746.58 895.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 854.88,750.00 C 861.28,743.60 868.14,736.74 870.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 885.12,750.00 C 878.72,756.40 871.86,763.26 870.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 930.00,775.20 C 919.02,764.22 908.22,753.42 904.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,724.80 C 940.98,735.78 951.78,746.58 955.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,750.00 Q 937.32,753.03 943.20,750.00 Q 937.32,746.97 930.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,750.00 Q 933.03,757.32 939.33,759.33 Q 937.32,753.03 930.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,750.00 Q 926.97,757.32 930.00,763.20 Q 933.03,757.32 930.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,750.00 Q 922.68,753.03 920.67,759.33 Q 926.97,757.32 930.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,750.00 Q 922.68,746.97 916.80,750.00 Q 922.68,753.03 930.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,750.00 Q 926.97,742.68 920.67,740.67 Q 922.68,746.97 930.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,750.00 Q 933.03,742.68 930.00,736.80 Q 926.97,742.68 930.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,750.00 Q 937.32,746.97 939.33,740.67 Q 933.03,742.68 930.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,750.00 Q 930.93,753.48 935.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,750.00 Q 926.52,750.93 924.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,750.00 Q 929.07,746.52 924.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,750.00 Q 933.48,749.07 935.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 914.88,750.00 C 921.28,743.60 928.14,736.74 930.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 945.12,750.00 C 938.72,756.40 931.86,763.26 930.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,724.80 C 1000.98,735.78 1011.78,746.58 1015.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,775.20 C 979.02,764.22 968.22,753.42 964.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 990.00,750.00 Q 997.32,753.03 1003.20,750.00 Q 997.32,746.97 990.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,750.00 Q 993.03,757.32 999.33,759.33 Q 997.32,753.03 990.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,750.00 Q 986.97,757.32 990.00,763.20 Q 993.03,757.32 990.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,750.00 Q 982.68,753.03 980.67,759.33 Q 986.97,757.32 990.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,750.00 Q 982.68,746.97 976.80,750.00 Q 982.68,753.03 990.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,750.00 Q 986.97,742.68 980.67,740.67 Q 982.68,746.97 990.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,750.00 Q 993.03,742.68 990.00,736.80 Q 986.97,742.68 990.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,750.00 Q 997.32,746.97 999.33,740.67 Q 993.03,742.68 990.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,750.00 Q 990.93,753.48 995.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,750.00 Q 986.52,750.93 984.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,750.00 Q 989.07,746.52 984.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,750.00 Q 993.48,749.07 995.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="990.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1005.12,750.00 C 998.72,756.40 991.86,763.26 990.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 974.88,750.00 C 981.28,743.60 988.14,736.74 990.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1075.20,750.00 C 1064.22,760.98 1053.42,771.78 1050.00,775.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1024.80,750.00 C 1035.78,739.02 1046.58,728.22 1050.00,724.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,765.12 C 1043.60,758.72 1036.74,751.86 1034.88,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,734.88 C 1056.40,741.28 1063.26,748.14 1065.12,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1110.00,724.80 C 1120.98,735.78 1131.78,746.58 1135.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,775.20 C 1099.02,764.22 1088.22,753.42 1084.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1125.12,750.00 C 1118.72,756.40 1111.86,763.26 1110.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1094.88,750.00 C 1101.28,743.60 1108.14,736.74 1110.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1170.00,775.20 C 1159.02,764.22 1148.22,753.42 1144.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,724.80 C 1180.98,735.78 1191.78,746.58 1195.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1154.88,750.00 C 1161.28,743.60 1168.14,736.74 1170.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1185.12,750.00 C 1178.72,756.40 1171.86,763.26 1170.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,724.80 C 1240.98,735.78 1251.78,746.58 1255.20,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,775.20 C 1219.02,764.22 1208.22,753.42 1204.80,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1245.12,750.00 C 1238.72,756.40 1231.86,763.26 1230.00,765.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1214.88,750.00 C 1221.28,743.60 1228.14,736.74 1230.00,734.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1315.20,750.00 C 1304.22,760.98 1293.42,771.78 1290.00,775.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1264.80,750.00 C 1275.78,739.02 1286.58,728.22 1290.00,724.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1290.00,750.00 Q 1297.32,753.03 1303.20,750.00 Q 1297.32,746.97 1290.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,750.00 Q 1293.03,757.32 1299.33,759.33 Q 1297.32,753.03 1290.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,750.00 Q 1286.97,757.32 1290.00,763.20 Q 1293.03,757.32 1290.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,750.00 Q 1282.68,753.03 1280.67,759.33 Q 1286.97,757.32 1290.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,750.00 Q 1282.68,746.97 1276.80,750.00 Q 1282.68,753.03 1290.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,750.00 Q 1286.97,742.68 1280.67,740.67 Q 1282.68,746.97 1290.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,750.00 Q 1293.03,742.68 1290.00,736.80 Q 1286.97,742.68 1290.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,750.00 Q 1297.32,746.97 1299.33,740.67 Q 1293.03,742.68 1290.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,750.00 Q 1290.93,753.48 1295.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,750.00 Q 1286.52,750.93 1284.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,750.00 Q 1289.07,746.52 1284.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,750.00 Q 1293.48,749.07 1295.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1290.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1290.00,765.12 C 1283.60,758.72 1276.74,751.86 1274.88,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,734.88 C 1296.40,741.28 1303.26,748.14 1305.12,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1375.20,750.00 C 1364.22,760.98 1353.42,771.78 1350.00,775.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1324.80,750.00 C 1335.78,739.02 1346.58,728.22 1350.00,724.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1350.00,750.00 Q 1357.32,753.03 1363.20,750.00 Q 1357.32,746.97 1350.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,750.00 Q 1353.03,757.32 1359.33,759.33 Q 1357.32,753.03 1350.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,750.00 Q 1346.97,757.32 1350.00,763.20 Q 1353.03,757.32 1350.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,750.00 Q 1342.68,753.03 1340.67,759.33 Q 1346.97,757.32 1350.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,750.00 Q 1342.68,746.97 1336.80,750.00 Q 1342.68,753.03 1350.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,750.00 Q 1346.97,742.68 1340.67,740.67 Q 1342.68,746.97 1350.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,750.00 Q 1353.03,742.68 1350.00,736.80 Q 1346.97,742.68 1350.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,750.00 Q 1357.32,746.97 1359.33,740.67 Q 1353.03,742.68 1350.00,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,750.00 Q 1350.93,753.48 1355.09,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,750.00 Q 1346.52,750.93 1344.91,755.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,750.00 Q 1349.07,746.52 1344.91,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,750.00 Q 1353.48,749.07 1355.09,744.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1350.0" cy="750.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1350.00,765.12 C 1343.60,758.72 1336.74,751.86 1334.88,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,734.88 C 1356.40,741.28 1363.26,748.14 1365.12,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,835.20 C 139.02,824.22 128.22,813.42 124.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,784.80 C 160.98,795.78 171.78,806.58 175.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 134.88,810.00 C 141.28,803.60 148.14,796.74 150.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 165.12,810.00 C 158.72,816.40 151.86,823.26 150.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 210.00,784.80 C 220.98,795.78 231.78,806.58 235.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,835.20 C 199.02,824.22 188.22,813.42 184.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 210.00,810.00 Q 217.32,813.03 223.20,810.00 Q 217.32,806.97 210.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,810.00 Q 213.03,817.32 219.33,819.33 Q 217.32,813.03 210.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,810.00 Q 206.97,817.32 210.00,823.20 Q 213.03,817.32 210.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,810.00 Q 202.68,813.03 200.67,819.33 Q 206.97,817.32 210.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,810.00 Q 202.68,806.97 196.80,810.00 Q 202.68,813.03 210.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,810.00 Q 206.97,802.68 200.67,800.67 Q 202.68,806.97 210.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,810.00 Q 213.03,802.68 210.00,796.80 Q 206.97,802.68 210.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,810.00 Q 217.32,806.97 219.33,800.67 Q 213.03,802.68 210.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,810.00 Q 210.93,813.48 215.09,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,810.00 Q 206.52,810.93 204.91,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,810.00 Q 209.07,806.52 204.91,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,810.00 Q 213.48,809.07 215.09,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="210.0" cy="810.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 225.12,810.00 C 218.72,816.40 211.86,823.26 210.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 194.88,810.00 C 201.28,803.60 208.14,796.74 210.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,784.80 C 280.98,795.78 291.78,806.58 295.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,835.20 C 259.02,824.22 248.22,813.42 244.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 285.12,810.00 C 278.72,816.40 271.86,823.26 270.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 254.88,810.00 C 261.28,803.60 268.14,796.74 270.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 330.00,835.20 C 319.02,824.22 308.22,813.42 304.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,784.80 C 340.98,795.78 351.78,806.58 355.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 314.88,810.00 C 321.28,803.60 328.14,796.74 330.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 345.12,810.00 C 338.72,816.40 331.86,823.26 330.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 390.00,784.80 C 400.98,795.78 411.78,806.58 415.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,835.20 C 379.02,824.22 368.22,813.42 364.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 390.00,810.00 Q 397.32,813.03 403.20,810.00 Q 397.32,806.97 390.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,810.00 Q 393.03,817.32 399.33,819.33 Q 397.32,813.03 390.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,810.00 Q 386.97,817.32 390.00,823.20 Q 393.03,817.32 390.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,810.00 Q 382.68,813.03 380.67,819.33 Q 386.97,817.32 390.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,810.00 Q 382.68,806.97 376.80,810.00 Q 382.68,813.03 390.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,810.00 Q 386.97,802.68 380.67,800.67 Q 382.68,806.97 390.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,810.00 Q 393.03,802.68 390.00,796.80 Q 386.97,802.68 390.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,810.00 Q 397.32,806.97 399.33,800.67 Q 393.03,802.68 390.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,810.00 Q 390.93,813.48 395.09,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,810.00 Q 386.52,810.93 384.91,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,810.00 Q 389.07,806.52 384.91,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,810.00 Q 393.48,809.07 395.09,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="390.0" cy="810.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 405.12,810.00 C 398.72,816.40 391.86,823.26 390.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 374.88,810.00 C 381.28,803.60 388.14,796.74 390.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 424.80,810.00 C 435.78,799.02 446.58,788.22 450.00,784.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 475.20,810.00 C 464.22,820.98 453.42,831.78 450.00,835.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 450.00,810.00 Q 457.32,813.03 463.20,810.00 Q 457.32,806.97 450.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,810.00 Q 453.03,817.32 459.33,819.33 Q 457.32,813.03 450.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,810.00 Q 446.97,817.32 450.00,823.20 Q 453.03,817.32 450.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,810.00 Q 442.68,813.03 440.67,819.33 Q 446.97,817.32 450.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,810.00 Q 442.68,806.97 436.80,810.00 Q 442.68,813.03 450.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,810.00 Q 446.97,802.68 440.67,800.67 Q 442.68,806.97 450.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,810.00 Q 453.03,802.68 450.00,796.80 Q 446.97,802.68 450.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,810.00 Q 457.32,806.97 459.33,800.67 Q 453.03,802.68 450.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,810.00 Q 450.93,813.48 455.09,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,810.00 Q 446.52,810.93 444.91,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,810.00 Q 449.07,806.52 444.91,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,810.00 Q 453.48,809.07 455.09,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="450.0" cy="810.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 450.00,794.88 C 456.40,801.28 463.26,808.14 465.12,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,825.12 C 443.60,818.72 436.74,811.86 434.88,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 484.80,810.00 C 495.78,799.02 506.58,788.22 510.00,784.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 535.20,810.00 C 524.22,820.98 513.42,831.78 510.00,835.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 510.00,794.88 C 516.40,801.28 523.26,808.14 525.12,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,825.12 C 503.60,818.72 496.74,811.86 494.88,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 570.00,835.20 C 559.02,824.22 548.22,813.42 544.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,784.80 C 580.98,795.78 591.78,806.58 595.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 554.88,810.00 C 561.28,803.60 568.14,796.74 570.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 585.12,810.00 C 578.72,816.40 571.86,823.26 570.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 655.20,810.00 C 644.22,820.98 633.42,831.78 630.00,835.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 604.80,810.00 C 615.78,799.02 626.58,788.22 630.00,784.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,825.12 C 623.60,818.72 616.74,811.86 614.88,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,794.88 C 636.40,801.28 643.26,808.14 645.12,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 690.00,784.80 C 700.98,795.78 711.78,806.58 715.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,835.20 C 679.02,824.22 668.22,813.42 664.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 690.00,810.00 Q 697.32,813.03 703.20,810.00 Q 697.32,806.97 690.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,810.00 Q 693.03,817.32 699.33,819.33 Q 697.32,813.03 690.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,810.00 Q 686.97,817.32 690.00,823.20 Q 693.03,817.32 690.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,810.00 Q 682.68,813.03 680.67,819.33 Q 686.97,817.32 690.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,810.00 Q 682.68,806.97 676.80,810.00 Q 682.68,813.03 690.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,810.00 Q 686.97,802.68 680.67,800.67 Q 682.68,806.97 690.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,810.00 Q 693.03,802.68 690.00,796.80 Q 686.97,802.68 690.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,810.00 Q 697.32,806.97 699.33,800.67 Q 693.03,802.68 690.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,810.00 Q 690.93,813.48 695.09,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,810.00 Q 686.52,810.93 684.91,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,810.00 Q 689.07,806.52 684.91,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,810.00 Q 693.48,809.07 695.09,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="690.0" cy="810.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 705.12,810.00 C 698.72,816.40 691.86,823.26 690.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 674.88,810.00 C 681.28,803.60 688.14,796.74 690.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 775.20,810.00 C 764.22,820.98 753.42,831.78 750.00,835.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 724.80,810.00 C 735.78,799.02 746.58,788.22 750.00,784.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,825.12 C 743.60,818.72 736.74,811.86 734.88,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,794.88 C 756.40,801.28 763.26,808.14 765.12,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 835.20,810.00 C 824.22,820.98 813.42,831.78 810.00,835.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 784.80,810.00 C 795.78,799.02 806.58,788.22 810.00,784.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,825.12 C 803.60,818.72 796.74,811.86 794.88,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,794.88 C 816.40,801.28 823.26,808.14 825.12,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 870.00,784.80 C 880.98,795.78 891.78,806.58 895.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,835.20 C 859.02,824.22 848.22,813.42 844.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,810.00 Q 877.32,813.03 883.20,810.00 Q 877.32,806.97 870.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,810.00 Q 873.03,817.32 879.33,819.33 Q 877.32,813.03 870.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,810.00 Q 866.97,817.32 870.00,823.20 Q 873.03,817.32 870.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,810.00 Q 862.68,813.03 860.67,819.33 Q 866.97,817.32 870.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,810.00 Q 862.68,806.97 856.80,810.00 Q 862.68,813.03 870.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,810.00 Q 866.97,802.68 860.67,800.67 Q 862.68,806.97 870.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,810.00 Q 873.03,802.68 870.00,796.80 Q 866.97,802.68 870.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,810.00 Q 877.32,806.97 879.33,800.67 Q 873.03,802.68 870.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,810.00 Q 870.93,813.48 875.09,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,810.00 Q 866.52,810.93 864.91,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,810.00 Q 869.07,806.52 864.91,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,810.00 Q 873.48,809.07 875.09,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="810.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 885.12,810.00 C 878.72,816.40 871.86,823.26 870.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 854.88,810.00 C 861.28,803.60 868.14,796.74 870.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 904.80,810.00 C 915.78,799.02 926.58,788.22 930.00,784.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 955.20,810.00 C 944.22,820.98 933.42,831.78 930.00,835.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,810.00 Q 937.32,813.03 943.20,810.00 Q 937.32,806.97 930.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,810.00 Q 933.03,817.32 939.33,819.33 Q 937.32,813.03 930.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,810.00 Q 926.97,817.32 930.00,823.20 Q 933.03,817.32 930.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,810.00 Q 922.68,813.03 920.67,819.33 Q 926.97,817.32 930.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,810.00 Q 922.68,806.97 916.80,810.00 Q 922.68,813.03 930.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,810.00 Q 926.97,802.68 920.67,800.67 Q 922.68,806.97 930.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,810.00 Q 933.03,802.68 930.00,796.80 Q 926.97,802.68 930.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,810.00 Q 937.32,806.97 939.33,800.67 Q 933.03,802.68 930.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,810.00 Q 930.93,813.48 935.09,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,810.00 Q 926.52,810.93 924.91,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,810.00 Q 929.07,806.52 924.91,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,810.00 Q 933.48,809.07 935.09,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="810.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 930.00,794.88 C 936.40,801.28 943.26,808.14 945.12,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,825.12 C 923.60,818.72 916.74,811.86 914.88,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 964.80,810.00 C 975.78,799.02 986.58,788.22 990.00,784.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1015.20,810.00 C 1004.22,820.98 993.42,831.78 990.00,835.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 990.00,794.88 C 996.40,801.28 1003.26,808.14 1005.12,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,825.12 C 983.60,818.72 976.74,811.86 974.88,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1050.00,835.20 C 1039.02,824.22 1028.22,813.42 1024.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,784.80 C 1060.98,795.78 1071.78,806.58 1075.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1034.88,810.00 C 1041.28,803.60 1048.14,796.74 1050.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1065.12,810.00 C 1058.72,816.40 1051.86,823.26 1050.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1110.00,784.80 C 1120.98,795.78 1131.78,806.58 1135.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,835.20 C 1099.02,824.22 1088.22,813.42 1084.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1110.00,810.00 Q 1117.32,813.03 1123.20,810.00 Q 1117.32,806.97 1110.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,810.00 Q 1113.03,817.32 1119.33,819.33 Q 1117.32,813.03 1110.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,810.00 Q 1106.97,817.32 1110.00,823.20 Q 1113.03,817.32 1110.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,810.00 Q 1102.68,813.03 1100.67,819.33 Q 1106.97,817.32 1110.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,810.00 Q 1102.68,806.97 1096.80,810.00 Q 1102.68,813.03 1110.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,810.00 Q 1106.97,802.68 1100.67,800.67 Q 1102.68,806.97 1110.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,810.00 Q 1113.03,802.68 1110.00,796.80 Q 1106.97,802.68 1110.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,810.00 Q 1117.32,806.97 1119.33,800.67 Q 1113.03,802.68 1110.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,810.00 Q 1110.93,813.48 1115.09,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,810.00 Q 1106.52,810.93 1104.91,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,810.00 Q 1109.07,806.52 1104.91,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,810.00 Q 1113.48,809.07 1115.09,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1110.0" cy="810.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1125.12,810.00 C 1118.72,816.40 1111.86,823.26 1110.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1094.88,810.00 C 1101.28,803.60 1108.14,796.74 1110.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1170.00,784.80 C 1180.98,795.78 1191.78,806.58 1195.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,835.20 C 1159.02,824.22 1148.22,813.42 1144.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1170.00,810.00 Q 1177.32,813.03 1183.20,810.00 Q 1177.32,806.97 1170.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,810.00 Q 1173.03,817.32 1179.33,819.33 Q 1177.32,813.03 1170.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,810.00 Q 1166.97,817.32 1170.00,823.20 Q 1173.03,817.32 1170.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,810.00 Q 1162.68,813.03 1160.67,819.33 Q 1166.97,817.32 1170.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,810.00 Q 1162.68,806.97 1156.80,810.00 Q 1162.68,813.03 1170.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,810.00 Q 1166.97,802.68 1160.67,800.67 Q 1162.68,806.97 1170.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,810.00 Q 1173.03,802.68 1170.00,796.80 Q 1166.97,802.68 1170.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,810.00 Q 1177.32,806.97 1179.33,800.67 Q 1173.03,802.68 1170.00,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,810.00 Q 1170.93,813.48 1175.09,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,810.00 Q 1166.52,810.93 1164.91,815.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,810.00 Q 1169.07,806.52 1164.91,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,810.00 Q 1173.48,809.07 1175.09,804.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1170.0" cy="810.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1185.12,810.00 C 1178.72,816.40 1171.86,823.26 1170.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1154.88,810.00 C 1161.28,803.60 1168.14,796.74 1170.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1255.20,810.00 C 1244.22,820.98 1233.42,831.78 1230.00,835.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1204.80,810.00 C 1215.78,799.02 1226.58,788.22 1230.00,784.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1230.00,825.12 C 1223.60,818.72 1216.74,811.86 1214.88,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,794.88 C 1236.40,801.28 1243.26,808.14 1245.12,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1315.20,810.00 C 1304.22,820.98 1293.42,831.78 1290.00,835.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1264.80,810.00 C 1275.78,799.02 1286.58,788.22 1290.00,784.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1290.00,825.12 C 1283.60,818.72 1276.74,811.86 1274.88,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,794.88 C 1296.40,801.28 1303.26,808.14 1305.12,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1350.00,835.20 C 1339.02,824.22 1328.22,813.42 1324.80,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,784.80 C 1360.98,795.78 1371.78,806.58 1375.20,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1334.88,810.00 C 1341.28,803.60 1348.14,796.74 1350.00,794.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1365.12,810.00 C 1358.72,816.40 1351.86,823.26 1350.00,825.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,844.80 C 160.98,855.78 171.78,866.58 175.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,895.20 C 139.02,884.22 128.22,873.42 124.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,870.00 Q 157.32,873.03 163.20,870.00 Q 157.32,866.97 150.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,870.00 Q 153.03,877.32 159.33,879.33 Q 157.32,873.03 150.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,870.00 Q 146.97,877.32 150.00,883.20 Q 153.03,877.32 150.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,870.00 Q 142.68,873.03 140.67,879.33 Q 146.97,877.32 150.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,870.00 Q 142.68,866.97 136.80,870.00 Q 142.68,873.03 150.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,870.00 Q 146.97,862.68 140.67,860.67 Q 142.68,866.97 150.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,870.00 Q 153.03,862.68 150.00,856.80 Q 146.97,862.68 150.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,870.00 Q 157.32,866.97 159.33,860.67 Q 153.03,862.68 150.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,870.00 Q 150.93,873.48 155.09,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,870.00 Q 146.52,870.93 144.91,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,870.00 Q 149.07,866.52 144.91,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,870.00 Q 153.48,869.07 155.09,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="870.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 165.12,870.00 C 158.72,876.40 151.86,883.26 150.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 134.88,870.00 C 141.28,863.60 148.14,856.74 150.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 184.80,870.00 C 195.78,859.02 206.58,848.22 210.00,844.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 235.20,870.00 C 224.22,880.98 213.42,891.78 210.00,895.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,854.88 C 216.40,861.28 223.26,868.14 225.12,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,885.12 C 203.60,878.72 196.74,871.86 194.88,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,895.20 C 259.02,884.22 248.22,873.42 244.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,844.80 C 280.98,855.78 291.78,866.58 295.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 254.88,870.00 C 261.28,863.60 268.14,856.74 270.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 285.12,870.00 C 278.72,876.40 271.86,883.26 270.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 330.00,844.80 C 340.98,855.78 351.78,866.58 355.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,895.20 C 319.02,884.22 308.22,873.42 304.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 345.12,870.00 C 338.72,876.40 331.86,883.26 330.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 314.88,870.00 C 321.28,863.60 328.14,856.74 330.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,870.00 C 375.78,859.02 386.58,848.22 390.00,844.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,870.00 C 404.22,880.98 393.42,891.78 390.00,895.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 390.00,870.00 Q 397.32,873.03 403.20,870.00 Q 397.32,866.97 390.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,870.00 Q 393.03,877.32 399.33,879.33 Q 397.32,873.03 390.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,870.00 Q 386.97,877.32 390.00,883.20 Q 393.03,877.32 390.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,870.00 Q 382.68,873.03 380.67,879.33 Q 386.97,877.32 390.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,870.00 Q 382.68,866.97 376.80,870.00 Q 382.68,873.03 390.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,870.00 Q 386.97,862.68 380.67,860.67 Q 382.68,866.97 390.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,870.00 Q 393.03,862.68 390.00,856.80 Q 386.97,862.68 390.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,870.00 Q 397.32,866.97 399.33,860.67 Q 393.03,862.68 390.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,870.00 Q 390.93,873.48 395.09,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,870.00 Q 386.52,870.93 384.91,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,870.00 Q 389.07,866.52 384.91,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,870.00 Q 393.48,869.07 395.09,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="390.0" cy="870.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 390.00,854.88 C 396.40,861.28 403.26,868.14 405.12,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,885.12 C 383.60,878.72 376.74,871.86 374.88,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 475.20,870.00 C 464.22,880.98 453.42,891.78 450.00,895.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 424.80,870.00 C 435.78,859.02 446.58,848.22 450.00,844.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 450.00,885.12 C 443.60,878.72 436.74,871.86 434.88,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,854.88 C 456.40,861.28 463.26,868.14 465.12,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,895.20 C 499.02,884.22 488.22,873.42 484.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,844.80 C 520.98,855.78 531.78,866.58 535.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 494.88,870.00 C 501.28,863.60 508.14,856.74 510.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 525.12,870.00 C 518.72,876.40 511.86,883.26 510.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 570.00,844.80 C 580.98,855.78 591.78,866.58 595.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,895.20 C 559.02,884.22 548.22,873.42 544.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 585.12,870.00 C 578.72,876.40 571.86,883.26 570.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 554.88,870.00 C 561.28,863.60 568.14,856.74 570.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,870.00 C 615.78,859.02 626.58,848.22 630.00,844.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,870.00 C 644.22,880.98 633.42,891.78 630.00,895.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,854.88 C 636.40,861.28 643.26,868.14 645.12,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,885.12 C 623.60,878.72 616.74,871.86 614.88,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 664.80,870.00 C 675.78,859.02 686.58,848.22 690.00,844.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 715.20,870.00 C 704.22,880.98 693.42,891.78 690.00,895.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 690.00,854.88 C 696.40,861.28 703.26,868.14 705.12,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,885.12 C 683.60,878.72 676.74,871.86 674.88,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 750.00,895.20 C 739.02,884.22 728.22,873.42 724.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,844.80 C 760.98,855.78 771.78,866.58 775.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 734.88,870.00 C 741.28,863.60 748.14,856.74 750.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 765.12,870.00 C 758.72,876.40 751.86,883.26 750.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 835.20,870.00 C 824.22,880.98 813.42,891.78 810.00,895.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 784.80,870.00 C 795.78,859.02 806.58,848.22 810.00,844.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,885.12 C 803.60,878.72 796.74,871.86 794.88,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,854.88 C 816.40,861.28 823.26,868.14 825.12,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 870.00,844.80 C 880.98,855.78 891.78,866.58 895.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,895.20 C 859.02,884.22 848.22,873.42 844.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,870.00 Q 877.32,873.03 883.20,870.00 Q 877.32,866.97 870.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,870.00 Q 873.03,877.32 879.33,879.33 Q 877.32,873.03 870.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,870.00 Q 866.97,877.32 870.00,883.20 Q 873.03,877.32 870.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,870.00 Q 862.68,873.03 860.67,879.33 Q 866.97,877.32 870.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,870.00 Q 862.68,866.97 856.80,870.00 Q 862.68,873.03 870.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,870.00 Q 866.97,862.68 860.67,860.67 Q 862.68,866.97 870.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,870.00 Q 873.03,862.68 870.00,856.80 Q 866.97,862.68 870.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,870.00 Q 877.32,866.97 879.33,860.67 Q 873.03,862.68 870.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,870.00 Q 870.93,873.48 875.09,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,870.00 Q 866.52,870.93 864.91,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,870.00 Q 869.07,866.52 864.91,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,870.00 Q 873.48,869.07 875.09,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="870.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 885.12,870.00 C 878.72,876.40 871.86,883.26 870.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 854.88,870.00 C 861.28,863.60 868.14,856.74 870.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 930.00,844.80 C 940.98,855.78 951.78,866.58 955.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,895.20 C 919.02,884.22 908.22,873.42 904.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 945.12,870.00 C 938.72,876.40 931.86,883.26 930.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 914.88,870.00 C 921.28,863.60 928.14,856.74 930.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,895.20 C 979.02,884.22 968.22,873.42 964.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,844.80 C 1000.98,855.78 1011.78,866.58 1015.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 974.88,870.00 C 981.28,863.60 988.14,856.74 990.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1005.12,870.00 C 998.72,876.40 991.86,883.26 990.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1050.00,844.80 C 1060.98,855.78 1071.78,866.58 1075.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,895.20 C 1039.02,884.22 1028.22,873.42 1024.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1050.00,870.00 Q 1057.32,873.03 1063.20,870.00 Q 1057.32,866.97 1050.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,870.00 Q 1053.03,877.32 1059.33,879.33 Q 1057.32,873.03 1050.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,870.00 Q 1046.97,877.32 1050.00,883.20 Q 1053.03,877.32 1050.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,870.00 Q 1042.68,873.03 1040.67,879.33 Q 1046.97,877.32 1050.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,870.00 Q 1042.68,866.97 1036.80,870.00 Q 1042.68,873.03 1050.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,870.00 Q 1046.97,862.68 1040.67,860.67 Q 1042.68,866.97 1050.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,870.00 Q 1053.03,862.68 1050.00,856.80 Q 1046.97,862.68 1050.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,870.00 Q 1057.32,866.97 1059.33,860.67 Q 1053.03,862.68 1050.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,870.00 Q 1050.93,873.48 1055.09,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,870.00 Q 1046.52,870.93 1044.91,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,870.00 Q 1049.07,866.52 1044.91,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,870.00 Q 1053.48,869.07 1055.09,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1050.0" cy="870.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1065.12,870.00 C 1058.72,876.40 1051.86,883.26 1050.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1034.88,870.00 C 1041.28,863.60 1048.14,856.74 1050.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1084.80,870.00 C 1095.78,859.02 1106.58,848.22 1110.00,844.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1135.20,870.00 C 1124.22,880.98 1113.42,891.78 1110.00,895.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1110.00,870.00 Q 1117.32,873.03 1123.20,870.00 Q 1117.32,866.97 1110.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,870.00 Q 1113.03,877.32 1119.33,879.33 Q 1117.32,873.03 1110.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,870.00 Q 1106.97,877.32 1110.00,883.20 Q 1113.03,877.32 1110.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,870.00 Q 1102.68,873.03 1100.67,879.33 Q 1106.97,877.32 1110.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,870.00 Q 1102.68,866.97 1096.80,870.00 Q 1102.68,873.03 1110.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,870.00 Q 1106.97,862.68 1100.67,860.67 Q 1102.68,866.97 1110.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,870.00 Q 1113.03,862.68 1110.00,856.80 Q 1106.97,862.68 1110.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,870.00 Q 1117.32,866.97 1119.33,860.67 Q 1113.03,862.68 1110.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,870.00 Q 1110.93,873.48 1115.09,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,870.00 Q 1106.52,870.93 1104.91,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,870.00 Q 1109.07,866.52 1104.91,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,870.00 Q 1113.48,869.07 1115.09,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1110.0" cy="870.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1110.00,854.88 C 1116.40,861.28 1123.26,868.14 1125.12,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,885.12 C 1103.60,878.72 1096.74,871.86 1094.88,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1144.80,870.00 C 1155.78,859.02 1166.58,848.22 1170.00,844.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1195.20,870.00 C 1184.22,880.98 1173.42,891.78 1170.00,895.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1170.00,854.88 C 1176.40,861.28 1183.26,868.14 1185.12,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,885.12 C 1163.60,878.72 1156.74,871.86 1154.88,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,895.20 C 1219.02,884.22 1208.22,873.42 1204.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,844.80 C 1240.98,855.78 1251.78,866.58 1255.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1214.88,870.00 C 1221.28,863.60 1228.14,856.74 1230.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1245.12,870.00 C 1238.72,876.40 1231.86,883.26 1230.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1315.20,870.00 C 1304.22,880.98 1293.42,891.78 1290.00,895.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1264.80,870.00 C 1275.78,859.02 1286.58,848.22 1290.00,844.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1290.00,885.12 C 1283.60,878.72 1276.74,871.86 1274.88,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,854.88 C 1296.40,861.28 1303.26,868.14 1305.12,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1350.00,844.80 C 1360.98,855.78 1371.78,866.58 1375.20,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,895.20 C 1339.02,884.22 1328.22,873.42 1324.80,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1350.00,870.00 Q 1357.32,873.03 1363.20,870.00 Q 1357.32,866.97 1350.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,870.00 Q 1353.03,877.32 1359.33,879.33 Q 1357.32,873.03 1350.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,870.00 Q 1346.97,877.32 1350.00,883.20 Q 1353.03,877.32 1350.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,870.00 Q 1342.68,873.03 1340.67,879.33 Q 1346.97,877.32 1350.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,870.00 Q 1342.68,866.97 1336.80,870.00 Q 1342.68,873.03 1350.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,870.00 Q 1346.97,862.68 1340.67,860.67 Q 1342.68,866.97 1350.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,870.00 Q 1353.03,862.68 1350.00,856.80 Q 1346.97,862.68 1350.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,870.00 Q 1357.32,866.97 1359.33,860.67 Q 1353.03,862.68 1350.00,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,870.00 Q 1350.93,873.48 1355.09,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,870.00 Q 1346.52,870.93 1344.91,875.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,870.00 Q 1349.07,866.52 1344.91,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,870.00 Q 1353.48,869.07 1355.09,864.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1350.0" cy="870.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1365.12,870.00 C 1358.72,876.40 1351.86,883.26 1350.00,885.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1334.88,870.00 C 1341.28,863.60 1348.14,856.74 1350.00,854.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,904.80 C 160.98,915.78 171.78,926.58 175.20,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,955.20 C 139.02,944.22 128.22,933.42 124.80,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,930.00 Q 157.32,933.03 163.20,930.00 Q 157.32,926.97 150.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,930.00 Q 153.03,937.32 159.33,939.33 Q 157.32,933.03 150.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,930.00 Q 146.97,937.32 150.00,943.20 Q 153.03,937.32 150.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,930.00 Q 142.68,933.03 140.67,939.33 Q 146.97,937.32 150.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,930.00 Q 142.68,926.97 136.80,930.00 Q 142.68,933.03 150.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,930.00 Q 146.97,922.68 140.67,920.67 Q 142.68,926.97 150.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,930.00 Q 153.03,922.68 150.00,916.80 Q 146.97,922.68 150.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,930.00 Q 157.32,926.97 159.33,920.67 Q 153.03,922.68 150.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,930.00 Q 150.93,933.48 155.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,930.00 Q 146.52,930.93 144.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,930.00 Q 149.07,926.52 144.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,930.00 Q 153.48,929.07 155.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 165.12,930.00 C 158.72,936.40 151.86,943.26 150.00,945.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 134.88,930.00 C 141.28,923.60 148.14,916.74 150.00,914.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 235.20,930.00 C 224.22,940.98 213.42,951.78 210.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 184.80,930.00 C 195.78,919.02 206.58,908.22 210.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,945.12 C 203.60,938.72 196.74,931.86 194.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,914.88 C 216.40,921.28 223.26,928.14 225.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,955.20 C 259.02,944.22 248.22,933.42 244.80,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,904.80 C 280.98,915.78 291.78,926.58 295.20,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 254.88,930.00 C 261.28,923.60 268.14,916.74 270.00,914.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 285.12,930.00 C 278.72,936.40 271.86,943.26 270.00,945.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 330.00,955.20 C 319.02,944.22 308.22,933.42 304.80,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,904.80 C 340.98,915.78 351.78,926.58 355.20,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 330.00,930.00 Q 337.32,933.03 343.20,930.00 Q 337.32,926.97 330.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,930.00 Q 333.03,937.32 339.33,939.33 Q 337.32,933.03 330.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,930.00 Q 326.97,937.32 330.00,943.20 Q 333.03,937.32 330.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,930.00 Q 322.68,933.03 320.67,939.33 Q 326.97,937.32 330.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,930.00 Q 322.68,926.97 316.80,930.00 Q 322.68,933.03 330.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,930.00 Q 326.97,922.68 320.67,920.67 Q 322.68,926.97 330.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,930.00 Q 333.03,922.68 330.00,916.80 Q 326.97,922.68 330.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,930.00 Q 337.32,926.97 339.33,920.67 Q 333.03,922.68 330.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,930.00 Q 330.93,933.48 335.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,930.00 Q 326.52,930.93 324.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,930.00 Q 329.07,926.52 324.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,930.00 Q 333.48,929.07 335.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="330.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 314.88,930.00 C 321.28,923.60 328.14,916.74 330.00,914.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 345.12,930.00 C 338.72,936.40 331.86,943.26 330.00,945.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,930.00 C 375.78,919.02 386.58,908.22 390.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,930.00 C 404.22,940.98 393.42,951.78 390.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 390.00,914.88 C 396.40,921.28 403.26,928.14 405.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,945.12 C 383.60,938.72 376.74,931.86 374.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 475.20,930.00 C 464.22,940.98 453.42,951.78 450.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 424.80,930.00 C 435.78,919.02 446.58,908.22 450.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 450.00,945.12 C 443.60,938.72 436.74,931.86 434.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,914.88 C 456.40,921.28 463.26,928.14 465.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,904.80 C 520.98,915.78 531.78,926.58 535.20,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,955.20 C 499.02,944.22 488.22,933.42 484.80,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 510.00,930.00 Q 517.32,933.03 523.20,930.00 Q 517.32,926.97 510.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,930.00 Q 513.03,937.32 519.33,939.33 Q 517.32,933.03 510.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,930.00 Q 506.97,937.32 510.00,943.20 Q 513.03,937.32 510.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,930.00 Q 502.68,933.03 500.67,939.33 Q 506.97,937.32 510.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,930.00 Q 502.68,926.97 496.80,930.00 Q 502.68,933.03 510.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,930.00 Q 506.97,922.68 500.67,920.67 Q 502.68,926.97 510.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,930.00 Q 513.03,922.68 510.00,916.80 Q 506.97,922.68 510.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,930.00 Q 517.32,926.97 519.33,920.67 Q 513.03,922.68 510.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 510.00,930.00 Q 510.93,933.48 515.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,930.00 Q 506.52,930.93 504.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,930.00 Q 509.07,926.52 504.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 510.00,930.00 Q 513.48,929.07 515.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="510.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 525.12,930.00 C 518.72,936.40 511.86,943.26 510.00,945.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 494.88,930.00 C 501.28,923.60 508.14,916.74 510.00,914.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,930.00 C 555.78,919.02 566.58,908.22 570.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,930.00 C 584.22,940.98 573.42,951.78 570.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 570.00,930.00 Q 577.32,933.03 583.20,930.00 Q 577.32,926.97 570.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,930.00 Q 573.03,937.32 579.33,939.33 Q 577.32,933.03 570.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,930.00 Q 566.97,937.32 570.00,943.20 Q 573.03,937.32 570.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,930.00 Q 562.68,933.03 560.67,939.33 Q 566.97,937.32 570.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,930.00 Q 562.68,926.97 556.80,930.00 Q 562.68,933.03 570.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,930.00 Q 566.97,922.68 560.67,920.67 Q 562.68,926.97 570.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,930.00 Q 573.03,922.68 570.00,916.80 Q 566.97,922.68 570.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,930.00 Q 577.32,926.97 579.33,920.67 Q 573.03,922.68 570.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,930.00 Q 570.93,933.48 575.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,930.00 Q 566.52,930.93 564.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,930.00 Q 569.07,926.52 564.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,930.00 Q 573.48,929.07 575.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="570.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 570.00,914.88 C 576.40,921.28 583.26,928.14 585.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,945.12 C 563.60,938.72 556.74,931.86 554.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,930.00 C 615.78,919.02 626.58,908.22 630.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,930.00 C 644.22,940.98 633.42,951.78 630.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 630.00,930.00 Q 637.32,933.03 643.20,930.00 Q 637.32,926.97 630.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,930.00 Q 633.03,937.32 639.33,939.33 Q 637.32,933.03 630.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,930.00 Q 626.97,937.32 630.00,943.20 Q 633.03,937.32 630.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,930.00 Q 622.68,933.03 620.67,939.33 Q 626.97,937.32 630.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,930.00 Q 622.68,926.97 616.80,930.00 Q 622.68,933.03 630.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,930.00 Q 626.97,922.68 620.67,920.67 Q 622.68,926.97 630.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,930.00 Q 633.03,922.68 630.00,916.80 Q 626.97,922.68 630.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,930.00 Q 637.32,926.97 639.33,920.67 Q 633.03,922.68 630.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,930.00 Q 630.93,933.48 635.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,930.00 Q 626.52,930.93 624.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,930.00 Q 629.07,926.52 624.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,930.00 Q 633.48,929.07 635.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="630.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 630.00,914.88 C 636.40,921.28 643.26,928.14 645.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,945.12 C 623.60,938.72 616.74,931.86 614.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 664.80,930.00 C 675.78,919.02 686.58,908.22 690.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 715.20,930.00 C 704.22,940.98 693.42,951.78 690.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 690.00,914.88 C 696.40,921.28 703.26,928.14 705.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,945.12 C 683.60,938.72 676.74,931.86 674.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 750.00,904.80 C 760.98,915.78 771.78,926.58 775.20,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,955.20 C 739.02,944.22 728.22,933.42 724.80,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 765.12,930.00 C 758.72,936.40 751.86,943.26 750.00,945.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 734.88,930.00 C 741.28,923.60 748.14,916.74 750.00,914.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 784.80,930.00 C 795.78,919.02 806.58,908.22 810.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 835.20,930.00 C 824.22,940.98 813.42,951.78 810.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,914.88 C 816.40,921.28 823.26,928.14 825.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,945.12 C 803.60,938.72 796.74,931.86 794.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 844.80,930.00 C 855.78,919.02 866.58,908.22 870.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 895.20,930.00 C 884.22,940.98 873.42,951.78 870.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,930.00 Q 877.32,933.03 883.20,930.00 Q 877.32,926.97 870.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,930.00 Q 873.03,937.32 879.33,939.33 Q 877.32,933.03 870.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,930.00 Q 866.97,937.32 870.00,943.20 Q 873.03,937.32 870.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,930.00 Q 862.68,933.03 860.67,939.33 Q 866.97,937.32 870.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,930.00 Q 862.68,926.97 856.80,930.00 Q 862.68,933.03 870.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,930.00 Q 866.97,922.68 860.67,920.67 Q 862.68,926.97 870.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,930.00 Q 873.03,922.68 870.00,916.80 Q 866.97,922.68 870.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,930.00 Q 877.32,926.97 879.33,920.67 Q 873.03,922.68 870.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,930.00 Q 870.93,933.48 875.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,930.00 Q 866.52,930.93 864.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,930.00 Q 869.07,926.52 864.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,930.00 Q 873.48,929.07 875.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 870.00,914.88 C 876.40,921.28 883.26,928.14 885.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,945.12 C 863.60,938.72 856.74,931.86 854.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 955.20,930.00 C 944.22,940.98 933.42,951.78 930.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 904.80,930.00 C 915.78,919.02 926.58,908.22 930.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,930.00 Q 937.32,933.03 943.20,930.00 Q 937.32,926.97 930.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,930.00 Q 933.03,937.32 939.33,939.33 Q 937.32,933.03 930.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,930.00 Q 926.97,937.32 930.00,943.20 Q 933.03,937.32 930.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,930.00 Q 922.68,933.03 920.67,939.33 Q 926.97,937.32 930.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,930.00 Q 922.68,926.97 916.80,930.00 Q 922.68,933.03 930.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,930.00 Q 926.97,922.68 920.67,920.67 Q 922.68,926.97 930.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,930.00 Q 933.03,922.68 930.00,916.80 Q 926.97,922.68 930.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,930.00 Q 937.32,926.97 939.33,920.67 Q 933.03,922.68 930.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,930.00 Q 930.93,933.48 935.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,930.00 Q 926.52,930.93 924.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,930.00 Q 929.07,926.52 924.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,930.00 Q 933.48,929.07 935.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 930.00,945.12 C 923.60,938.72 916.74,931.86 914.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,914.88 C 936.40,921.28 943.26,928.14 945.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,904.80 C 1000.98,915.78 1011.78,926.58 1015.20,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,955.20 C 979.02,944.22 968.22,933.42 964.80,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 990.00,930.00 Q 997.32,933.03 1003.20,930.00 Q 997.32,926.97 990.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,930.00 Q 993.03,937.32 999.33,939.33 Q 997.32,933.03 990.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,930.00 Q 986.97,937.32 990.00,943.20 Q 993.03,937.32 990.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,930.00 Q 982.68,933.03 980.67,939.33 Q 986.97,937.32 990.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,930.00 Q 982.68,926.97 976.80,930.00 Q 982.68,933.03 990.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,930.00 Q 986.97,922.68 980.67,920.67 Q 982.68,926.97 990.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,930.00 Q 993.03,922.68 990.00,916.80 Q 986.97,922.68 990.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,930.00 Q 997.32,926.97 999.33,920.67 Q 993.03,922.68 990.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,930.00 Q 990.93,933.48 995.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,930.00 Q 986.52,930.93 984.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,930.00 Q 989.07,926.52 984.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,930.00 Q 993.48,929.07 995.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="990.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1005.12,930.00 C 998.72,936.40 991.86,943.26 990.00,945.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 974.88,930.00 C 981.28,923.60 988.14,916.74 990.00,914.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,930.00 C 1035.78,919.02 1046.58,908.22 1050.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,930.00 C 1064.22,940.98 1053.42,951.78 1050.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1050.00,930.00 Q 1057.32,933.03 1063.20,930.00 Q 1057.32,926.97 1050.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,930.00 Q 1053.03,937.32 1059.33,939.33 Q 1057.32,933.03 1050.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,930.00 Q 1046.97,937.32 1050.00,943.20 Q 1053.03,937.32 1050.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,930.00 Q 1042.68,933.03 1040.67,939.33 Q 1046.97,937.32 1050.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,930.00 Q 1042.68,926.97 1036.80,930.00 Q 1042.68,933.03 1050.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,930.00 Q 1046.97,922.68 1040.67,920.67 Q 1042.68,926.97 1050.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,930.00 Q 1053.03,922.68 1050.00,916.80 Q 1046.97,922.68 1050.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,930.00 Q 1057.32,926.97 1059.33,920.67 Q 1053.03,922.68 1050.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,930.00 Q 1050.93,933.48 1055.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,930.00 Q 1046.52,930.93 1044.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,930.00 Q 1049.07,926.52 1044.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,930.00 Q 1053.48,929.07 1055.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1050.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1050.00,914.88 C 1056.40,921.28 1063.26,928.14 1065.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,945.12 C 1043.60,938.72 1036.74,931.86 1034.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1135.20,930.00 C 1124.22,940.98 1113.42,951.78 1110.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1084.80,930.00 C 1095.78,919.02 1106.58,908.22 1110.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1110.00,945.12 C 1103.60,938.72 1096.74,931.86 1094.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,914.88 C 1116.40,921.28 1123.26,928.14 1125.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1170.00,955.20 C 1159.02,944.22 1148.22,933.42 1144.80,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,904.80 C 1180.98,915.78 1191.78,926.58 1195.20,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1154.88,930.00 C 1161.28,923.60 1168.14,916.74 1170.00,914.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1185.12,930.00 C 1178.72,936.40 1171.86,943.26 1170.00,945.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,955.20 C 1219.02,944.22 1208.22,933.42 1204.80,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,904.80 C 1240.98,915.78 1251.78,926.58 1255.20,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1230.00,930.00 Q 1237.32,933.03 1243.20,930.00 Q 1237.32,926.97 1230.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,930.00 Q 1233.03,937.32 1239.33,939.33 Q 1237.32,933.03 1230.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,930.00 Q 1226.97,937.32 1230.00,943.20 Q 1233.03,937.32 1230.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,930.00 Q 1222.68,933.03 1220.67,939.33 Q 1226.97,937.32 1230.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,930.00 Q 1222.68,926.97 1216.80,930.00 Q 1222.68,933.03 1230.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,930.00 Q 1226.97,922.68 1220.67,920.67 Q 1222.68,926.97 1230.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,930.00 Q 1233.03,922.68 1230.00,916.80 Q 1226.97,922.68 1230.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,930.00 Q 1237.32,926.97 1239.33,920.67 Q 1233.03,922.68 1230.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,930.00 Q 1230.93,933.48 1235.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,930.00 Q 1226.52,930.93 1224.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,930.00 Q 1229.07,926.52 1224.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,930.00 Q 1233.48,929.07 1235.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1230.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1214.88,930.00 C 1221.28,923.60 1228.14,916.74 1230.00,914.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1245.12,930.00 C 1238.72,936.40 1231.86,943.26 1230.00,945.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1290.00,904.80 C 1300.98,915.78 1311.78,926.58 1315.20,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,955.20 C 1279.02,944.22 1268.22,933.42 1264.80,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1290.00,930.00 Q 1297.32,933.03 1303.20,930.00 Q 1297.32,926.97 1290.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,930.00 Q 1293.03,937.32 1299.33,939.33 Q 1297.32,933.03 1290.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,930.00 Q 1286.97,937.32 1290.00,943.20 Q 1293.03,937.32 1290.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,930.00 Q 1282.68,933.03 1280.67,939.33 Q 1286.97,937.32 1290.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,930.00 Q 1282.68,926.97 1276.80,930.00 Q 1282.68,933.03 1290.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,930.00 Q 1286.97,922.68 1280.67,920.67 Q 1282.68,926.97 1290.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,930.00 Q 1293.03,922.68 1290.00,916.80 Q 1286.97,922.68 1290.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,930.00 Q 1297.32,926.97 1299.33,920.67 Q 1293.03,922.68 1290.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,930.00 Q 1290.93,933.48 1295.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,930.00 Q 1286.52,930.93 1284.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,930.00 Q 1289.07,926.52 1284.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,930.00 Q 1293.48,929.07 1295.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1290.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1305.12,930.00 C 1298.72,936.40 1291.86,943.26 1290.00,945.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1274.88,930.00 C 1281.28,923.60 1288.14,916.74 1290.00,914.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1375.20,930.00 C 1364.22,940.98 1353.42,951.78 1350.00,955.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1324.80,930.00 C 1335.78,919.02 1346.58,908.22 1350.00,904.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1350.00,930.00 Q 1357.32,933.03 1363.20,930.00 Q 1357.32,926.97 1350.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,930.00 Q 1353.03,937.32 1359.33,939.33 Q 1357.32,933.03 1350.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,930.00 Q 1346.97,937.32 1350.00,943.20 Q 1353.03,937.32 1350.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,930.00 Q 1342.68,933.03 1340.67,939.33 Q 1346.97,937.32 1350.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,930.00 Q 1342.68,926.97 1336.80,930.00 Q 1342.68,933.03 1350.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,930.00 Q 1346.97,922.68 1340.67,920.67 Q 1342.68,926.97 1350.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,930.00 Q 1353.03,922.68 1350.00,916.80 Q 1346.97,922.68 1350.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,930.00 Q 1357.32,926.97 1359.33,920.67 Q 1353.03,922.68 1350.00,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,930.00 Q 1350.93,933.48 1355.09,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,930.00 Q 1346.52,930.93 1344.91,935.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,930.00 Q 1349.07,926.52 1344.91,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,930.00 Q 1353.48,929.07 1355.09,924.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1350.0" cy="930.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1350.00,945.12 C 1343.60,938.72 1336.74,931.86 1334.88,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,914.88 C 1356.40,921.28 1363.26,928.14 1365.12,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 175.20,990.00 C 164.22,1000.98 153.42,1011.78 150.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 124.80,990.00 C 135.78,979.02 146.58,968.22 150.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 150.00,1005.12 C 143.60,998.72 136.74,991.86 134.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,974.88 C 156.40,981.28 163.26,988.14 165.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 235.20,990.00 C 224.22,1000.98 213.42,1011.78 210.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 184.80,990.00 C 195.78,979.02 206.58,968.22 210.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 210.00,990.00 Q 217.32,993.03 223.20,990.00 Q 217.32,986.97 210.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,990.00 Q 213.03,997.32 219.33,999.33 Q 217.32,993.03 210.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,990.00 Q 206.97,997.32 210.00,1003.20 Q 213.03,997.32 210.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,990.00 Q 202.68,993.03 200.67,999.33 Q 206.97,997.32 210.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,990.00 Q 202.68,986.97 196.80,990.00 Q 202.68,993.03 210.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,990.00 Q 206.97,982.68 200.67,980.67 Q 202.68,986.97 210.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,990.00 Q 213.03,982.68 210.00,976.80 Q 206.97,982.68 210.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,990.00 Q 217.32,986.97 219.33,980.67 Q 213.03,982.68 210.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,990.00 Q 210.93,993.48 215.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,990.00 Q 206.52,990.93 204.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,990.00 Q 209.07,986.52 204.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,990.00 Q 213.48,989.07 215.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="210.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 210.00,1005.12 C 203.60,998.72 196.74,991.86 194.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,974.88 C 216.40,981.28 223.26,988.14 225.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,964.80 C 280.98,975.78 291.78,986.58 295.20,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,1015.20 C 259.02,1004.22 248.22,993.42 244.80,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 270.00,990.00 Q 277.32,993.03 283.20,990.00 Q 277.32,986.97 270.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,990.00 Q 273.03,997.32 279.33,999.33 Q 277.32,993.03 270.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,990.00 Q 266.97,997.32 270.00,1003.20 Q 273.03,997.32 270.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,990.00 Q 262.68,993.03 260.67,999.33 Q 266.97,997.32 270.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,990.00 Q 262.68,986.97 256.80,990.00 Q 262.68,993.03 270.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,990.00 Q 266.97,982.68 260.67,980.67 Q 262.68,986.97 270.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,990.00 Q 273.03,982.68 270.00,976.80 Q 266.97,982.68 270.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,990.00 Q 277.32,986.97 279.33,980.67 Q 273.03,982.68 270.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,990.00 Q 270.93,993.48 275.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,990.00 Q 266.52,990.93 264.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,990.00 Q 269.07,986.52 264.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,990.00 Q 273.48,989.07 275.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="270.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 285.12,990.00 C 278.72,996.40 271.86,1003.26 270.00,1005.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 254.88,990.00 C 261.28,983.60 268.14,976.74 270.00,974.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,990.00 C 315.78,979.02 326.58,968.22 330.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,990.00 C 344.22,1000.98 333.42,1011.78 330.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 330.00,990.00 Q 337.32,993.03 343.20,990.00 Q 337.32,986.97 330.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,990.00 Q 333.03,997.32 339.33,999.33 Q 337.32,993.03 330.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,990.00 Q 326.97,997.32 330.00,1003.20 Q 333.03,997.32 330.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,990.00 Q 322.68,993.03 320.67,999.33 Q 326.97,997.32 330.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,990.00 Q 322.68,986.97 316.80,990.00 Q 322.68,993.03 330.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,990.00 Q 326.97,982.68 320.67,980.67 Q 322.68,986.97 330.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,990.00 Q 333.03,982.68 330.00,976.80 Q 326.97,982.68 330.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,990.00 Q 337.32,986.97 339.33,980.67 Q 333.03,982.68 330.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 330.00,990.00 Q 330.93,993.48 335.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,990.00 Q 326.52,990.93 324.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,990.00 Q 329.07,986.52 324.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 330.00,990.00 Q 333.48,989.07 335.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="330.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 330.00,974.88 C 336.40,981.28 343.26,988.14 345.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,1005.12 C 323.60,998.72 316.74,991.86 314.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 415.20,990.00 C 404.22,1000.98 393.42,1011.78 390.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 364.80,990.00 C 375.78,979.02 386.58,968.22 390.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 390.00,1005.12 C 383.60,998.72 376.74,991.86 374.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,974.88 C 396.40,981.28 403.26,988.14 405.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 450.00,1015.20 C 439.02,1004.22 428.22,993.42 424.80,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,964.80 C 460.98,975.78 471.78,986.58 475.20,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 434.88,990.00 C 441.28,983.60 448.14,976.74 450.00,974.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 465.12,990.00 C 458.72,996.40 451.86,1003.26 450.00,1005.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 510.00,964.80 C 520.98,975.78 531.78,986.58 535.20,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,1015.20 C 499.02,1004.22 488.22,993.42 484.80,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 525.12,990.00 C 518.72,996.40 511.86,1003.26 510.00,1005.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 494.88,990.00 C 501.28,983.60 508.14,976.74 510.00,974.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 595.20,990.00 C 584.22,1000.98 573.42,1011.78 570.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 544.80,990.00 C 555.78,979.02 566.58,968.22 570.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 570.00,990.00 Q 577.32,993.03 583.20,990.00 Q 577.32,986.97 570.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,990.00 Q 573.03,997.32 579.33,999.33 Q 577.32,993.03 570.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,990.00 Q 566.97,997.32 570.00,1003.20 Q 573.03,997.32 570.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,990.00 Q 562.68,993.03 560.67,999.33 Q 566.97,997.32 570.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,990.00 Q 562.68,986.97 556.80,990.00 Q 562.68,993.03 570.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,990.00 Q 566.97,982.68 560.67,980.67 Q 562.68,986.97 570.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,990.00 Q 573.03,982.68 570.00,976.80 Q 566.97,982.68 570.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,990.00 Q 577.32,986.97 579.33,980.67 Q 573.03,982.68 570.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 570.00,990.00 Q 570.93,993.48 575.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,990.00 Q 566.52,990.93 564.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,990.00 Q 569.07,986.52 564.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 570.00,990.00 Q 573.48,989.07 575.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="570.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 570.00,1005.12 C 563.60,998.72 556.74,991.86 554.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,974.88 C 576.40,981.28 583.26,988.14 585.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 630.00,1015.20 C 619.02,1004.22 608.22,993.42 604.80,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,964.80 C 640.98,975.78 651.78,986.58 655.20,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 614.88,990.00 C 621.28,983.60 628.14,976.74 630.00,974.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 645.12,990.00 C 638.72,996.40 631.86,1003.26 630.00,1005.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 690.00,1015.20 C 679.02,1004.22 668.22,993.42 664.80,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,964.80 C 700.98,975.78 711.78,986.58 715.20,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 690.00,990.00 Q 697.32,993.03 703.20,990.00 Q 697.32,986.97 690.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,990.00 Q 693.03,997.32 699.33,999.33 Q 697.32,993.03 690.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,990.00 Q 686.97,997.32 690.00,1003.20 Q 693.03,997.32 690.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,990.00 Q 682.68,993.03 680.67,999.33 Q 686.97,997.32 690.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,990.00 Q 682.68,986.97 676.80,990.00 Q 682.68,993.03 690.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,990.00 Q 686.97,982.68 680.67,980.67 Q 682.68,986.97 690.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,990.00 Q 693.03,982.68 690.00,976.80 Q 686.97,982.68 690.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,990.00 Q 697.32,986.97 699.33,980.67 Q 693.03,982.68 690.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,990.00 Q 690.93,993.48 695.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,990.00 Q 686.52,990.93 684.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,990.00 Q 689.07,986.52 684.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,990.00 Q 693.48,989.07 695.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="690.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 674.88,990.00 C 681.28,983.60 688.14,976.74 690.00,974.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 705.12,990.00 C 698.72,996.40 691.86,1003.26 690.00,1005.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 750.00,964.80 C 760.98,975.78 771.78,986.58 775.20,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,1015.20 C 739.02,1004.22 728.22,993.42 724.80,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 750.00,990.00 Q 757.32,993.03 763.20,990.00 Q 757.32,986.97 750.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,990.00 Q 753.03,997.32 759.33,999.33 Q 757.32,993.03 750.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,990.00 Q 746.97,997.32 750.00,1003.20 Q 753.03,997.32 750.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,990.00 Q 742.68,993.03 740.67,999.33 Q 746.97,997.32 750.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,990.00 Q 742.68,986.97 736.80,990.00 Q 742.68,993.03 750.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,990.00 Q 746.97,982.68 740.67,980.67 Q 742.68,986.97 750.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,990.00 Q 753.03,982.68 750.00,976.80 Q 746.97,982.68 750.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,990.00 Q 757.32,986.97 759.33,980.67 Q 753.03,982.68 750.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,990.00 Q 750.93,993.48 755.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,990.00 Q 746.52,990.93 744.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,990.00 Q 749.07,986.52 744.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,990.00 Q 753.48,989.07 755.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="750.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 765.12,990.00 C 758.72,996.40 751.86,1003.26 750.00,1005.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 734.88,990.00 C 741.28,983.60 748.14,976.74 750.00,974.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 835.20,990.00 C 824.22,1000.98 813.42,1011.78 810.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 784.80,990.00 C 795.78,979.02 806.58,968.22 810.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,1005.12 C 803.60,998.72 796.74,991.86 794.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,974.88 C 816.40,981.28 823.26,988.14 825.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 895.20,990.00 C 884.22,1000.98 873.42,1011.78 870.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 844.80,990.00 C 855.78,979.02 866.58,968.22 870.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 870.00,1005.12 C 863.60,998.72 856.74,991.86 854.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,974.88 C 876.40,981.28 883.26,988.14 885.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 930.00,1015.20 C 919.02,1004.22 908.22,993.42 904.80,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,964.80 C 940.98,975.78 951.78,986.58 955.20,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 914.88,990.00 C 921.28,983.60 928.14,976.74 930.00,974.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 945.12,990.00 C 938.72,996.40 931.86,1003.26 930.00,1005.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,964.80 C 1000.98,975.78 1011.78,986.58 1015.20,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,1015.20 C 979.02,1004.22 968.22,993.42 964.80,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 990.00,990.00 Q 997.32,993.03 1003.20,990.00 Q 997.32,986.97 990.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,990.00 Q 993.03,997.32 999.33,999.33 Q 997.32,993.03 990.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,990.00 Q 986.97,997.32 990.00,1003.20 Q 993.03,997.32 990.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,990.00 Q 982.68,993.03 980.67,999.33 Q 986.97,997.32 990.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,990.00 Q 982.68,986.97 976.80,990.00 Q 982.68,993.03 990.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,990.00 Q 986.97,982.68 980.67,980.67 Q 982.68,986.97 990.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,990.00 Q 993.03,982.68 990.00,976.80 Q 986.97,982.68 990.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,990.00 Q 997.32,986.97 999.33,980.67 Q 993.03,982.68 990.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,990.00 Q 990.93,993.48 995.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,990.00 Q 986.52,990.93 984.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,990.00 Q 989.07,986.52 984.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,990.00 Q 993.48,989.07 995.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="990.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1005.12,990.00 C 998.72,996.40 991.86,1003.26 990.00,1005.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 974.88,990.00 C 981.28,983.60 988.14,976.74 990.00,974.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,990.00 C 1035.78,979.02 1046.58,968.22 1050.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,990.00 C 1064.22,1000.98 1053.42,1011.78 1050.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1050.00,990.00 Q 1057.32,993.03 1063.20,990.00 Q 1057.32,986.97 1050.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,990.00 Q 1053.03,997.32 1059.33,999.33 Q 1057.32,993.03 1050.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,990.00 Q 1046.97,997.32 1050.00,1003.20 Q 1053.03,997.32 1050.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,990.00 Q 1042.68,993.03 1040.67,999.33 Q 1046.97,997.32 1050.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,990.00 Q 1042.68,986.97 1036.80,990.00 Q 1042.68,993.03 1050.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,990.00 Q 1046.97,982.68 1040.67,980.67 Q 1042.68,986.97 1050.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,990.00 Q 1053.03,982.68 1050.00,976.80 Q 1046.97,982.68 1050.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,990.00 Q 1057.32,986.97 1059.33,980.67 Q 1053.03,982.68 1050.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,990.00 Q 1050.93,993.48 1055.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,990.00 Q 1046.52,990.93 1044.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,990.00 Q 1049.07,986.52 1044.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,990.00 Q 1053.48,989.07 1055.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1050.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1050.00,974.88 C 1056.40,981.28 1063.26,988.14 1065.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,1005.12 C 1043.60,998.72 1036.74,991.86 1034.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1135.20,990.00 C 1124.22,1000.98 1113.42,1011.78 1110.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1084.80,990.00 C 1095.78,979.02 1106.58,968.22 1110.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1110.00,1005.12 C 1103.60,998.72 1096.74,991.86 1094.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,974.88 C 1116.40,981.28 1123.26,988.14 1125.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1195.20,990.00 C 1184.22,1000.98 1173.42,1011.78 1170.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1144.80,990.00 C 1155.78,979.02 1166.58,968.22 1170.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1170.00,990.00 Q 1177.32,993.03 1183.20,990.00 Q 1177.32,986.97 1170.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,990.00 Q 1173.03,997.32 1179.33,999.33 Q 1177.32,993.03 1170.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,990.00 Q 1166.97,997.32 1170.00,1003.20 Q 1173.03,997.32 1170.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,990.00 Q 1162.68,993.03 1160.67,999.33 Q 1166.97,997.32 1170.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,990.00 Q 1162.68,986.97 1156.80,990.00 Q 1162.68,993.03 1170.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,990.00 Q 1166.97,982.68 1160.67,980.67 Q 1162.68,986.97 1170.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,990.00 Q 1173.03,982.68 1170.00,976.80 Q 1166.97,982.68 1170.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,990.00 Q 1177.32,986.97 1179.33,980.67 Q 1173.03,982.68 1170.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,990.00 Q 1170.93,993.48 1175.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,990.00 Q 1166.52,990.93 1164.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,990.00 Q 1169.07,986.52 1164.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,990.00 Q 1173.48,989.07 1175.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1170.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1170.00,1005.12 C 1163.60,998.72 1156.74,991.86 1154.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,974.88 C 1176.40,981.28 1183.26,988.14 1185.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1230.00,964.80 C 1240.98,975.78 1251.78,986.58 1255.20,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,1015.20 C 1219.02,1004.22 1208.22,993.42 1204.80,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1230.00,990.00 Q 1237.32,993.03 1243.20,990.00 Q 1237.32,986.97 1230.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,990.00 Q 1233.03,997.32 1239.33,999.33 Q 1237.32,993.03 1230.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,990.00 Q 1226.97,997.32 1230.00,1003.20 Q 1233.03,997.32 1230.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,990.00 Q 1222.68,993.03 1220.67,999.33 Q 1226.97,997.32 1230.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,990.00 Q 1222.68,986.97 1216.80,990.00 Q 1222.68,993.03 1230.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,990.00 Q 1226.97,982.68 1220.67,980.67 Q 1222.68,986.97 1230.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,990.00 Q 1233.03,982.68 1230.00,976.80 Q 1226.97,982.68 1230.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,990.00 Q 1237.32,986.97 1239.33,980.67 Q 1233.03,982.68 1230.00,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,990.00 Q 1230.93,993.48 1235.09,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,990.00 Q 1226.52,990.93 1224.91,995.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,990.00 Q 1229.07,986.52 1224.91,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,990.00 Q 1233.48,989.07 1235.09,984.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1230.0" cy="990.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1245.12,990.00 C 1238.72,996.40 1231.86,1003.26 1230.00,1005.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1214.88,990.00 C 1221.28,983.60 1228.14,976.74 1230.00,974.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1315.20,990.00 C 1304.22,1000.98 1293.42,1011.78 1290.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1264.80,990.00 C 1275.78,979.02 1286.58,968.22 1290.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1290.00,1005.12 C 1283.60,998.72 1276.74,991.86 1274.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,974.88 C 1296.40,981.28 1303.26,988.14 1305.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1375.20,990.00 C 1364.22,1000.98 1353.42,1011.78 1350.00,1015.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1324.80,990.00 C 1335.78,979.02 1346.58,968.22 1350.00,964.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,1005.12 C 1343.60,998.72 1336.74,991.86 1334.88,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,974.88 C 1356.40,981.28 1363.26,988.14 1365.12,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,1075.20 C 139.02,1064.22 128.22,1053.42 124.80,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,1024.80 C 160.98,1035.78 171.78,1046.58 175.20,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,1050.00 Q 157.32,1053.03 163.20,1050.00 Q 157.32,1046.97 150.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1050.00 Q 153.03,1057.32 159.33,1059.33 Q 157.32,1053.03 150.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1050.00 Q 146.97,1057.32 150.00,1063.20 Q 153.03,1057.32 150.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1050.00 Q 142.68,1053.03 140.67,1059.33 Q 146.97,1057.32 150.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1050.00 Q 142.68,1046.97 136.80,1050.00 Q 142.68,1053.03 150.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1050.00 Q 146.97,1042.68 140.67,1040.67 Q 142.68,1046.97 150.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1050.00 Q 153.03,1042.68 150.00,1036.80 Q 146.97,1042.68 150.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1050.00 Q 157.32,1046.97 159.33,1040.67 Q 153.03,1042.68 150.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1050.00 Q 150.93,1053.48 155.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,1050.00 Q 146.52,1050.93 144.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,1050.00 Q 149.07,1046.52 144.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,1050.00 Q 153.48,1049.07 155.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 134.88,1050.00 C 141.28,1043.60 148.14,1036.74 150.00,1034.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 165.12,1050.00 C 158.72,1056.40 151.86,1063.26 150.00,1065.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 210.00,1024.80 C 220.98,1035.78 231.78,1046.58 235.20,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,1075.20 C 199.02,1064.22 188.22,1053.42 184.80,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 210.00,1050.00 Q 217.32,1053.03 223.20,1050.00 Q 217.32,1046.97 210.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1050.00 Q 213.03,1057.32 219.33,1059.33 Q 217.32,1053.03 210.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1050.00 Q 206.97,1057.32 210.00,1063.20 Q 213.03,1057.32 210.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1050.00 Q 202.68,1053.03 200.67,1059.33 Q 206.97,1057.32 210.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1050.00 Q 202.68,1046.97 196.80,1050.00 Q 202.68,1053.03 210.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1050.00 Q 206.97,1042.68 200.67,1040.67 Q 202.68,1046.97 210.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1050.00 Q 213.03,1042.68 210.00,1036.80 Q 206.97,1042.68 210.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1050.00 Q 217.32,1046.97 219.33,1040.67 Q 213.03,1042.68 210.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1050.00 Q 210.93,1053.48 215.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,1050.00 Q 206.52,1050.93 204.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,1050.00 Q 209.07,1046.52 204.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,1050.00 Q 213.48,1049.07 215.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="210.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 225.12,1050.00 C 218.72,1056.40 211.86,1063.26 210.00,1065.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 194.88,1050.00 C 201.28,1043.60 208.14,1036.74 210.00,1034.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 244.80,1050.00 C 255.78,1039.02 266.58,1028.22 270.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 295.20,1050.00 C 284.22,1060.98 273.42,1071.78 270.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 270.00,1050.00 Q 277.32,1053.03 283.20,1050.00 Q 277.32,1046.97 270.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,1050.00 Q 273.03,1057.32 279.33,1059.33 Q 277.32,1053.03 270.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,1050.00 Q 266.97,1057.32 270.00,1063.20 Q 273.03,1057.32 270.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,1050.00 Q 262.68,1053.03 260.67,1059.33 Q 266.97,1057.32 270.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,1050.00 Q 262.68,1046.97 256.80,1050.00 Q 262.68,1053.03 270.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,1050.00 Q 266.97,1042.68 260.67,1040.67 Q 262.68,1046.97 270.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,1050.00 Q 273.03,1042.68 270.00,1036.80 Q 266.97,1042.68 270.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,1050.00 Q 277.32,1046.97 279.33,1040.67 Q 273.03,1042.68 270.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 270.00,1050.00 Q 270.93,1053.48 275.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,1050.00 Q 266.52,1050.93 264.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,1050.00 Q 269.07,1046.52 264.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 270.00,1050.00 Q 273.48,1049.07 275.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="270.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 270.00,1034.88 C 276.40,1041.28 283.26,1048.14 285.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,1065.12 C 263.60,1058.72 256.74,1051.86 254.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 330.00,1075.20 C 319.02,1064.22 308.22,1053.42 304.80,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,1024.80 C 340.98,1035.78 351.78,1046.58 355.20,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 314.88,1050.00 C 321.28,1043.60 328.14,1036.74 330.00,1034.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 345.12,1050.00 C 338.72,1056.40 331.86,1063.26 330.00,1065.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 390.00,1024.80 C 400.98,1035.78 411.78,1046.58 415.20,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,1075.20 C 379.02,1064.22 368.22,1053.42 364.80,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 405.12,1050.00 C 398.72,1056.40 391.86,1063.26 390.00,1065.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 374.88,1050.00 C 381.28,1043.60 388.14,1036.74 390.00,1034.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 424.80,1050.00 C 435.78,1039.02 446.58,1028.22 450.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 475.20,1050.00 C 464.22,1060.98 453.42,1071.78 450.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 450.00,1050.00 Q 457.32,1053.03 463.20,1050.00 Q 457.32,1046.97 450.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,1050.00 Q 453.03,1057.32 459.33,1059.33 Q 457.32,1053.03 450.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,1050.00 Q 446.97,1057.32 450.00,1063.20 Q 453.03,1057.32 450.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,1050.00 Q 442.68,1053.03 440.67,1059.33 Q 446.97,1057.32 450.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,1050.00 Q 442.68,1046.97 436.80,1050.00 Q 442.68,1053.03 450.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,1050.00 Q 446.97,1042.68 440.67,1040.67 Q 442.68,1046.97 450.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,1050.00 Q 453.03,1042.68 450.00,1036.80 Q 446.97,1042.68 450.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,1050.00 Q 457.32,1046.97 459.33,1040.67 Q 453.03,1042.68 450.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 450.00,1050.00 Q 450.93,1053.48 455.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,1050.00 Q 446.52,1050.93 444.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,1050.00 Q 449.07,1046.52 444.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 450.00,1050.00 Q 453.48,1049.07 455.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="450.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 450.00,1034.88 C 456.40,1041.28 463.26,1048.14 465.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,1065.12 C 443.60,1058.72 436.74,1051.86 434.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 484.80,1050.00 C 495.78,1039.02 506.58,1028.22 510.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 535.20,1050.00 C 524.22,1060.98 513.42,1071.78 510.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 510.00,1034.88 C 516.40,1041.28 523.26,1048.14 525.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,1065.12 C 503.60,1058.72 496.74,1051.86 494.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,1050.00 C 555.78,1039.02 566.58,1028.22 570.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,1050.00 C 584.22,1060.98 573.42,1071.78 570.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 570.00,1034.88 C 576.40,1041.28 583.26,1048.14 585.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,1065.12 C 563.60,1058.72 556.74,1051.86 554.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 630.00,1075.20 C 619.02,1064.22 608.22,1053.42 604.80,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,1024.80 C 640.98,1035.78 651.78,1046.58 655.20,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 614.88,1050.00 C 621.28,1043.60 628.14,1036.74 630.00,1034.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 645.12,1050.00 C 638.72,1056.40 631.86,1063.26 630.00,1065.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 664.80,1050.00 C 675.78,1039.02 686.58,1028.22 690.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 715.20,1050.00 C 704.22,1060.98 693.42,1071.78 690.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 690.00,1050.00 Q 697.32,1053.03 703.20,1050.00 Q 697.32,1046.97 690.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,1050.00 Q 693.03,1057.32 699.33,1059.33 Q 697.32,1053.03 690.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,1050.00 Q 686.97,1057.32 690.00,1063.20 Q 693.03,1057.32 690.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,1050.00 Q 682.68,1053.03 680.67,1059.33 Q 686.97,1057.32 690.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,1050.00 Q 682.68,1046.97 676.80,1050.00 Q 682.68,1053.03 690.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,1050.00 Q 686.97,1042.68 680.67,1040.67 Q 682.68,1046.97 690.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,1050.00 Q 693.03,1042.68 690.00,1036.80 Q 686.97,1042.68 690.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,1050.00 Q 697.32,1046.97 699.33,1040.67 Q 693.03,1042.68 690.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 690.00,1050.00 Q 690.93,1053.48 695.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,1050.00 Q 686.52,1050.93 684.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,1050.00 Q 689.07,1046.52 684.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 690.00,1050.00 Q 693.48,1049.07 695.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="690.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 690.00,1034.88 C 696.40,1041.28 703.26,1048.14 705.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,1065.12 C 683.60,1058.72 676.74,1051.86 674.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 724.80,1050.00 C 735.78,1039.02 746.58,1028.22 750.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 775.20,1050.00 C 764.22,1060.98 753.42,1071.78 750.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 750.00,1050.00 Q 757.32,1053.03 763.20,1050.00 Q 757.32,1046.97 750.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,1050.00 Q 753.03,1057.32 759.33,1059.33 Q 757.32,1053.03 750.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,1050.00 Q 746.97,1057.32 750.00,1063.20 Q 753.03,1057.32 750.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,1050.00 Q 742.68,1053.03 740.67,1059.33 Q 746.97,1057.32 750.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,1050.00 Q 742.68,1046.97 736.80,1050.00 Q 742.68,1053.03 750.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,1050.00 Q 746.97,1042.68 740.67,1040.67 Q 742.68,1046.97 750.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,1050.00 Q 753.03,1042.68 750.00,1036.80 Q 746.97,1042.68 750.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,1050.00 Q 757.32,1046.97 759.33,1040.67 Q 753.03,1042.68 750.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 750.00,1050.00 Q 750.93,1053.48 755.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,1050.00 Q 746.52,1050.93 744.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,1050.00 Q 749.07,1046.52 744.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 750.00,1050.00 Q 753.48,1049.07 755.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="750.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 750.00,1034.88 C 756.40,1041.28 763.26,1048.14 765.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,1065.12 C 743.60,1058.72 736.74,1051.86 734.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 835.20,1050.00 C 824.22,1060.98 813.42,1071.78 810.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 784.80,1050.00 C 795.78,1039.02 806.58,1028.22 810.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,1065.12 C 803.60,1058.72 796.74,1051.86 794.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,1034.88 C 816.40,1041.28 823.26,1048.14 825.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 870.00,1024.80 C 880.98,1035.78 891.78,1046.58 895.20,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,1075.20 C 859.02,1064.22 848.22,1053.42 844.80,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 885.12,1050.00 C 878.72,1056.40 871.86,1063.26 870.00,1065.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 854.88,1050.00 C 861.28,1043.60 868.14,1036.74 870.00,1034.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 904.80,1050.00 C 915.78,1039.02 926.58,1028.22 930.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 955.20,1050.00 C 944.22,1060.98 933.42,1071.78 930.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 930.00,1050.00 Q 937.32,1053.03 943.20,1050.00 Q 937.32,1046.97 930.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,1050.00 Q 933.03,1057.32 939.33,1059.33 Q 937.32,1053.03 930.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,1050.00 Q 926.97,1057.32 930.00,1063.20 Q 933.03,1057.32 930.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,1050.00 Q 922.68,1053.03 920.67,1059.33 Q 926.97,1057.32 930.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,1050.00 Q 922.68,1046.97 916.80,1050.00 Q 922.68,1053.03 930.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,1050.00 Q 926.97,1042.68 920.67,1040.67 Q 922.68,1046.97 930.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,1050.00 Q 933.03,1042.68 930.00,1036.80 Q 926.97,1042.68 930.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,1050.00 Q 937.32,1046.97 939.33,1040.67 Q 933.03,1042.68 930.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 930.00,1050.00 Q 930.93,1053.48 935.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,1050.00 Q 926.52,1050.93 924.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,1050.00 Q 929.07,1046.52 924.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 930.00,1050.00 Q 933.48,1049.07 935.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="930.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 930.00,1034.88 C 936.40,1041.28 943.26,1048.14 945.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,1065.12 C 923.60,1058.72 916.74,1051.86 914.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 964.80,1050.00 C 975.78,1039.02 986.58,1028.22 990.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1015.20,1050.00 C 1004.22,1060.98 993.42,1071.78 990.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 990.00,1034.88 C 996.40,1041.28 1003.26,1048.14 1005.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,1065.12 C 983.60,1058.72 976.74,1051.86 974.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,1050.00 C 1035.78,1039.02 1046.58,1028.22 1050.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,1050.00 C 1064.22,1060.98 1053.42,1071.78 1050.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,1034.88 C 1056.40,1041.28 1063.26,1048.14 1065.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,1065.12 C 1043.60,1058.72 1036.74,1051.86 1034.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1110.00,1075.20 C 1099.02,1064.22 1088.22,1053.42 1084.80,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,1024.80 C 1120.98,1035.78 1131.78,1046.58 1135.20,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1110.00,1050.00 Q 1117.32,1053.03 1123.20,1050.00 Q 1117.32,1046.97 1110.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,1050.00 Q 1113.03,1057.32 1119.33,1059.33 Q 1117.32,1053.03 1110.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,1050.00 Q 1106.97,1057.32 1110.00,1063.20 Q 1113.03,1057.32 1110.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,1050.00 Q 1102.68,1053.03 1100.67,1059.33 Q 1106.97,1057.32 1110.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,1050.00 Q 1102.68,1046.97 1096.80,1050.00 Q 1102.68,1053.03 1110.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,1050.00 Q 1106.97,1042.68 1100.67,1040.67 Q 1102.68,1046.97 1110.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,1050.00 Q 1113.03,1042.68 1110.00,1036.80 Q 1106.97,1042.68 1110.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,1050.00 Q 1117.32,1046.97 1119.33,1040.67 Q 1113.03,1042.68 1110.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1110.00,1050.00 Q 1110.93,1053.48 1115.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,1050.00 Q 1106.52,1050.93 1104.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,1050.00 Q 1109.07,1046.52 1104.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1110.00,1050.00 Q 1113.48,1049.07 1115.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1110.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1094.88,1050.00 C 1101.28,1043.60 1108.14,1036.74 1110.00,1034.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1125.12,1050.00 C 1118.72,1056.40 1111.86,1063.26 1110.00,1065.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1144.80,1050.00 C 1155.78,1039.02 1166.58,1028.22 1170.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1195.20,1050.00 C 1184.22,1060.98 1173.42,1071.78 1170.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1170.00,1050.00 Q 1177.32,1053.03 1183.20,1050.00 Q 1177.32,1046.97 1170.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,1050.00 Q 1173.03,1057.32 1179.33,1059.33 Q 1177.32,1053.03 1170.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,1050.00 Q 1166.97,1057.32 1170.00,1063.20 Q 1173.03,1057.32 1170.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,1050.00 Q 1162.68,1053.03 1160.67,1059.33 Q 1166.97,1057.32 1170.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,1050.00 Q 1162.68,1046.97 1156.80,1050.00 Q 1162.68,1053.03 1170.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,1050.00 Q 1166.97,1042.68 1160.67,1040.67 Q 1162.68,1046.97 1170.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,1050.00 Q 1173.03,1042.68 1170.00,1036.80 Q 1166.97,1042.68 1170.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,1050.00 Q 1177.32,1046.97 1179.33,1040.67 Q 1173.03,1042.68 1170.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1170.00,1050.00 Q 1170.93,1053.48 1175.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,1050.00 Q 1166.52,1050.93 1164.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,1050.00 Q 1169.07,1046.52 1164.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1170.00,1050.00 Q 1173.48,1049.07 1175.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1170.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1170.00,1034.88 C 1176.40,1041.28 1183.26,1048.14 1185.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,1065.12 C 1163.60,1058.72 1156.74,1051.86 1154.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1204.80,1050.00 C 1215.78,1039.02 1226.58,1028.22 1230.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1255.20,1050.00 C 1244.22,1060.98 1233.42,1071.78 1230.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1230.00,1050.00 Q 1237.32,1053.03 1243.20,1050.00 Q 1237.32,1046.97 1230.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1050.00 Q 1233.03,1057.32 1239.33,1059.33 Q 1237.32,1053.03 1230.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1050.00 Q 1226.97,1057.32 1230.00,1063.20 Q 1233.03,1057.32 1230.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1050.00 Q 1222.68,1053.03 1220.67,1059.33 Q 1226.97,1057.32 1230.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1050.00 Q 1222.68,1046.97 1216.80,1050.00 Q 1222.68,1053.03 1230.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1050.00 Q 1226.97,1042.68 1220.67,1040.67 Q 1222.68,1046.97 1230.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1050.00 Q 1233.03,1042.68 1230.00,1036.80 Q 1226.97,1042.68 1230.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1050.00 Q 1237.32,1046.97 1239.33,1040.67 Q 1233.03,1042.68 1230.00,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1050.00 Q 1230.93,1053.48 1235.09,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,1050.00 Q 1226.52,1050.93 1224.91,1055.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,1050.00 Q 1229.07,1046.52 1224.91,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,1050.00 Q 1233.48,1049.07 1235.09,1044.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1230.0" cy="1050.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1230.00,1034.88 C 1236.40,1041.28 1243.26,1048.14 1245.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,1065.12 C 1223.60,1058.72 1216.74,1051.86 1214.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1290.00,1075.20 C 1279.02,1064.22 1268.22,1053.42 1264.80,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,1024.80 C 1300.98,1035.78 1311.78,1046.58 1315.20,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1274.88,1050.00 C 1281.28,1043.60 1288.14,1036.74 1290.00,1034.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1305.12,1050.00 C 1298.72,1056.40 1291.86,1063.26 1290.00,1065.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1375.20,1050.00 C 1364.22,1060.98 1353.42,1071.78 1350.00,1075.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1324.80,1050.00 C 1335.78,1039.02 1346.58,1028.22 1350.00,1024.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,1065.12 C 1343.60,1058.72 1336.74,1051.86 1334.88,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,1034.88 C 1356.40,1041.28 1363.26,1048.14 1365.12,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 150.00,1084.80 C 160.98,1095.78 171.78,1106.58 175.20,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,1135.20 C 139.02,1124.22 128.22,1113.42 124.80,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 150.00,1110.00 Q 157.32,1113.03 163.20,1110.00 Q 157.32,1106.97 150.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1110.00 Q 153.03,1117.32 159.33,1119.33 Q 157.32,1113.03 150.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1110.00 Q 146.97,1117.32 150.00,1123.20 Q 153.03,1117.32 150.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1110.00 Q 142.68,1113.03 140.67,1119.33 Q 146.97,1117.32 150.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1110.00 Q 142.68,1106.97 136.80,1110.00 Q 142.68,1113.03 150.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1110.00 Q 146.97,1102.68 140.67,1100.67 Q 142.68,1106.97 150.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1110.00 Q 153.03,1102.68 150.00,1096.80 Q 146.97,1102.68 150.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1110.00 Q 157.32,1106.97 159.33,1100.67 Q 153.03,1102.68 150.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 150.00,1110.00 Q 150.93,1113.48 155.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,1110.00 Q 146.52,1110.93 144.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,1110.00 Q 149.07,1106.52 144.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 150.00,1110.00 Q 153.48,1109.07 155.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="150.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 165.12,1110.00 C 158.72,1116.40 151.86,1123.26 150.00,1125.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 134.88,1110.00 C 141.28,1103.60 148.14,1096.74 150.00,1094.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 184.80,1110.00 C 195.78,1099.02 206.58,1088.22 210.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 235.20,1110.00 C 224.22,1120.98 213.42,1131.78 210.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 210.00,1110.00 Q 217.32,1113.03 223.20,1110.00 Q 217.32,1106.97 210.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1110.00 Q 213.03,1117.32 219.33,1119.33 Q 217.32,1113.03 210.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1110.00 Q 206.97,1117.32 210.00,1123.20 Q 213.03,1117.32 210.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1110.00 Q 202.68,1113.03 200.67,1119.33 Q 206.97,1117.32 210.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1110.00 Q 202.68,1106.97 196.80,1110.00 Q 202.68,1113.03 210.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1110.00 Q 206.97,1102.68 200.67,1100.67 Q 202.68,1106.97 210.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1110.00 Q 213.03,1102.68 210.00,1096.80 Q 206.97,1102.68 210.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1110.00 Q 217.32,1106.97 219.33,1100.67 Q 213.03,1102.68 210.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 210.00,1110.00 Q 210.93,1113.48 215.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,1110.00 Q 206.52,1110.93 204.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,1110.00 Q 209.07,1106.52 204.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 210.00,1110.00 Q 213.48,1109.07 215.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="210.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 210.00,1094.88 C 216.40,1101.28 223.26,1108.14 225.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,1125.12 C 203.60,1118.72 196.74,1111.86 194.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 270.00,1135.20 C 259.02,1124.22 248.22,1113.42 244.80,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,1084.80 C 280.98,1095.78 291.78,1106.58 295.20,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 254.88,1110.00 C 261.28,1103.60 268.14,1096.74 270.00,1094.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 285.12,1110.00 C 278.72,1116.40 271.86,1123.26 270.00,1125.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 330.00,1135.20 C 319.02,1124.22 308.22,1113.42 304.80,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,1084.80 C 340.98,1095.78 351.78,1106.58 355.20,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 314.88,1110.00 C 321.28,1103.60 328.14,1096.74 330.00,1094.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 345.12,1110.00 C 338.72,1116.40 331.86,1123.26 330.00,1125.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,1110.00 C 375.78,1099.02 386.58,1088.22 390.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,1110.00 C 404.22,1120.98 393.42,1131.78 390.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 390.00,1110.00 Q 397.32,1113.03 403.20,1110.00 Q 397.32,1106.97 390.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,1110.00 Q 393.03,1117.32 399.33,1119.33 Q 397.32,1113.03 390.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,1110.00 Q 386.97,1117.32 390.00,1123.20 Q 393.03,1117.32 390.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,1110.00 Q 382.68,1113.03 380.67,1119.33 Q 386.97,1117.32 390.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,1110.00 Q 382.68,1106.97 376.80,1110.00 Q 382.68,1113.03 390.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,1110.00 Q 386.97,1102.68 380.67,1100.67 Q 382.68,1106.97 390.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,1110.00 Q 393.03,1102.68 390.00,1096.80 Q 386.97,1102.68 390.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,1110.00 Q 397.32,1106.97 399.33,1100.67 Q 393.03,1102.68 390.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 390.00,1110.00 Q 390.93,1113.48 395.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,1110.00 Q 386.52,1110.93 384.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,1110.00 Q 389.07,1106.52 384.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 390.00,1110.00 Q 393.48,1109.07 395.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="390.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 390.00,1094.88 C 396.40,1101.28 403.26,1108.14 405.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,1125.12 C 383.60,1118.72 376.74,1111.86 374.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 424.80,1110.00 C 435.78,1099.02 446.58,1088.22 450.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 475.20,1110.00 C 464.22,1120.98 453.42,1131.78 450.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 450.00,1094.88 C 456.40,1101.28 463.26,1108.14 465.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,1125.12 C 443.60,1118.72 436.74,1111.86 434.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 535.20,1110.00 C 524.22,1120.98 513.42,1131.78 510.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 484.80,1110.00 C 495.78,1099.02 506.58,1088.22 510.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 510.00,1125.12 C 503.60,1118.72 496.74,1111.86 494.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,1094.88 C 516.40,1101.28 523.26,1108.14 525.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,1110.00 C 555.78,1099.02 566.58,1088.22 570.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,1110.00 C 584.22,1120.98 573.42,1131.78 570.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 570.00,1094.88 C 576.40,1101.28 583.26,1108.14 585.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,1125.12 C 563.60,1118.72 556.74,1111.86 554.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 630.00,1084.80 C 640.98,1095.78 651.78,1106.58 655.20,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,1135.20 C 619.02,1124.22 608.22,1113.42 604.80,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 630.00,1110.00 Q 637.32,1113.03 643.20,1110.00 Q 637.32,1106.97 630.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,1110.00 Q 633.03,1117.32 639.33,1119.33 Q 637.32,1113.03 630.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,1110.00 Q 626.97,1117.32 630.00,1123.20 Q 633.03,1117.32 630.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,1110.00 Q 622.68,1113.03 620.67,1119.33 Q 626.97,1117.32 630.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,1110.00 Q 622.68,1106.97 616.80,1110.00 Q 622.68,1113.03 630.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,1110.00 Q 626.97,1102.68 620.67,1100.67 Q 622.68,1106.97 630.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,1110.00 Q 633.03,1102.68 630.00,1096.80 Q 626.97,1102.68 630.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,1110.00 Q 637.32,1106.97 639.33,1100.67 Q 633.03,1102.68 630.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 630.00,1110.00 Q 630.93,1113.48 635.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,1110.00 Q 626.52,1110.93 624.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,1110.00 Q 629.07,1106.52 624.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 630.00,1110.00 Q 633.48,1109.07 635.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="630.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 645.12,1110.00 C 638.72,1116.40 631.86,1123.26 630.00,1125.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 614.88,1110.00 C 621.28,1103.60 628.14,1096.74 630.00,1094.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 715.20,1110.00 C 704.22,1120.98 693.42,1131.78 690.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 664.80,1110.00 C 675.78,1099.02 686.58,1088.22 690.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 690.00,1125.12 C 683.60,1118.72 676.74,1111.86 674.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,1094.88 C 696.40,1101.28 703.26,1108.14 705.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 775.20,1110.00 C 764.22,1120.98 753.42,1131.78 750.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 724.80,1110.00 C 735.78,1099.02 746.58,1088.22 750.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,1125.12 C 743.60,1118.72 736.74,1111.86 734.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,1094.88 C 756.40,1101.28 763.26,1108.14 765.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 835.20,1110.00 C 824.22,1120.98 813.42,1131.78 810.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 784.80,1110.00 C 795.78,1099.02 806.58,1088.22 810.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 810.00,1110.00 Q 817.32,1113.03 823.20,1110.00 Q 817.32,1106.97 810.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,1110.00 Q 813.03,1117.32 819.33,1119.33 Q 817.32,1113.03 810.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,1110.00 Q 806.97,1117.32 810.00,1123.20 Q 813.03,1117.32 810.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,1110.00 Q 802.68,1113.03 800.67,1119.33 Q 806.97,1117.32 810.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,1110.00 Q 802.68,1106.97 796.80,1110.00 Q 802.68,1113.03 810.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,1110.00 Q 806.97,1102.68 800.67,1100.67 Q 802.68,1106.97 810.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,1110.00 Q 813.03,1102.68 810.00,1096.80 Q 806.97,1102.68 810.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,1110.00 Q 817.32,1106.97 819.33,1100.67 Q 813.03,1102.68 810.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 810.00,1110.00 Q 810.93,1113.48 815.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,1110.00 Q 806.52,1110.93 804.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,1110.00 Q 809.07,1106.52 804.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 810.00,1110.00 Q 813.48,1109.07 815.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="810.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 810.00,1125.12 C 803.60,1118.72 796.74,1111.86 794.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,1094.88 C 816.40,1101.28 823.26,1108.14 825.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 870.00,1084.80 C 880.98,1095.78 891.78,1106.58 895.20,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,1135.20 C 859.02,1124.22 848.22,1113.42 844.80,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 870.00,1110.00 Q 877.32,1113.03 883.20,1110.00 Q 877.32,1106.97 870.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,1110.00 Q 873.03,1117.32 879.33,1119.33 Q 877.32,1113.03 870.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,1110.00 Q 866.97,1117.32 870.00,1123.20 Q 873.03,1117.32 870.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,1110.00 Q 862.68,1113.03 860.67,1119.33 Q 866.97,1117.32 870.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,1110.00 Q 862.68,1106.97 856.80,1110.00 Q 862.68,1113.03 870.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,1110.00 Q 866.97,1102.68 860.67,1100.67 Q 862.68,1106.97 870.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,1110.00 Q 873.03,1102.68 870.00,1096.80 Q 866.97,1102.68 870.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,1110.00 Q 877.32,1106.97 879.33,1100.67 Q 873.03,1102.68 870.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 870.00,1110.00 Q 870.93,1113.48 875.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,1110.00 Q 866.52,1110.93 864.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,1110.00 Q 869.07,1106.52 864.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 870.00,1110.00 Q 873.48,1109.07 875.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="870.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 885.12,1110.00 C 878.72,1116.40 871.86,1123.26 870.00,1125.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 854.88,1110.00 C 861.28,1103.60 868.14,1096.74 870.00,1094.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 955.20,1110.00 C 944.22,1120.98 933.42,1131.78 930.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 904.80,1110.00 C 915.78,1099.02 926.58,1088.22 930.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 930.00,1125.12 C 923.60,1118.72 916.74,1111.86 914.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,1094.88 C 936.40,1101.28 943.26,1108.14 945.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 990.00,1084.80 C 1000.98,1095.78 1011.78,1106.58 1015.20,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,1135.20 C 979.02,1124.22 968.22,1113.42 964.80,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 990.00,1110.00 Q 997.32,1113.03 1003.20,1110.00 Q 997.32,1106.97 990.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,1110.00 Q 993.03,1117.32 999.33,1119.33 Q 997.32,1113.03 990.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,1110.00 Q 986.97,1117.32 990.00,1123.20 Q 993.03,1117.32 990.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,1110.00 Q 982.68,1113.03 980.67,1119.33 Q 986.97,1117.32 990.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,1110.00 Q 982.68,1106.97 976.80,1110.00 Q 982.68,1113.03 990.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,1110.00 Q 986.97,1102.68 980.67,1100.67 Q 982.68,1106.97 990.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,1110.00 Q 993.03,1102.68 990.00,1096.80 Q 986.97,1102.68 990.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,1110.00 Q 997.32,1106.97 999.33,1100.67 Q 993.03,1102.68 990.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 990.00,1110.00 Q 990.93,1113.48 995.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,1110.00 Q 986.52,1110.93 984.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,1110.00 Q 989.07,1106.52 984.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 990.00,1110.00 Q 993.48,1109.07 995.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="990.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1005.12,1110.00 C 998.72,1116.40 991.86,1123.26 990.00,1125.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 974.88,1110.00 C 981.28,1103.60 988.14,1096.74 990.00,1094.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1075.20,1110.00 C 1064.22,1120.98 1053.42,1131.78 1050.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1024.80,1110.00 C 1035.78,1099.02 1046.58,1088.22 1050.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1050.00,1110.00 Q 1057.32,1113.03 1063.20,1110.00 Q 1057.32,1106.97 1050.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,1110.00 Q 1053.03,1117.32 1059.33,1119.33 Q 1057.32,1113.03 1050.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,1110.00 Q 1046.97,1117.32 1050.00,1123.20 Q 1053.03,1117.32 1050.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,1110.00 Q 1042.68,1113.03 1040.67,1119.33 Q 1046.97,1117.32 1050.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,1110.00 Q 1042.68,1106.97 1036.80,1110.00 Q 1042.68,1113.03 1050.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,1110.00 Q 1046.97,1102.68 1040.67,1100.67 Q 1042.68,1106.97 1050.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,1110.00 Q 1053.03,1102.68 1050.00,1096.80 Q 1046.97,1102.68 1050.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,1110.00 Q 1057.32,1106.97 1059.33,1100.67 Q 1053.03,1102.68 1050.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1050.00,1110.00 Q 1050.93,1113.48 1055.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,1110.00 Q 1046.52,1110.93 1044.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,1110.00 Q 1049.07,1106.52 1044.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1050.00,1110.00 Q 1053.48,1109.07 1055.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1050.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1050.00,1125.12 C 1043.60,1118.72 1036.74,1111.86 1034.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,1094.88 C 1056.40,1101.28 1063.26,1108.14 1065.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1110.00,1084.80 C 1120.98,1095.78 1131.78,1106.58 1135.20,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,1135.20 C 1099.02,1124.22 1088.22,1113.42 1084.80,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1125.12,1110.00 C 1118.72,1116.40 1111.86,1123.26 1110.00,1125.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1094.88,1110.00 C 1101.28,1103.60 1108.14,1096.74 1110.00,1094.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1195.20,1110.00 C 1184.22,1120.98 1173.42,1131.78 1170.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1144.80,1110.00 C 1155.78,1099.02 1166.58,1088.22 1170.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1170.00,1125.12 C 1163.60,1118.72 1156.74,1111.86 1154.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,1094.88 C 1176.40,1101.28 1183.26,1108.14 1185.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1255.20,1110.00 C 1244.22,1120.98 1233.42,1131.78 1230.00,1135.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1204.80,1110.00 C 1215.78,1099.02 1226.58,1088.22 1230.00,1084.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1230.00,1110.00 Q 1237.32,1113.03 1243.20,1110.00 Q 1237.32,1106.97 1230.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1110.00 Q 1233.03,1117.32 1239.33,1119.33 Q 1237.32,1113.03 1230.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1110.00 Q 1226.97,1117.32 1230.00,1123.20 Q 1233.03,1117.32 1230.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1110.00 Q 1222.68,1113.03 1220.67,1119.33 Q 1226.97,1117.32 1230.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1110.00 Q 1222.68,1106.97 1216.80,1110.00 Q 1222.68,1113.03 1230.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1110.00 Q 1226.97,1102.68 1220.67,1100.67 Q 1222.68,1106.97 1230.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1110.00 Q 1233.03,1102.68 1230.00,1096.80 Q 1226.97,1102.68 1230.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1110.00 Q 1237.32,1106.97 1239.33,1100.67 Q 1233.03,1102.68 1230.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1230.00,1110.00 Q 1230.93,1113.48 1235.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,1110.00 Q 1226.52,1110.93 1224.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,1110.00 Q 1229.07,1106.52 1224.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1230.00,1110.00 Q 1233.48,1109.07 1235.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1230.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1230.00,1125.12 C 1223.60,1118.72 1216.74,1111.86 1214.88,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,1094.88 C 1236.40,1101.28 1243.26,1108.14 1245.12,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1290.00,1135.20 C 1279.02,1124.22 1268.22,1113.42 1264.80,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,1084.80 C 1300.98,1095.78 1311.78,1106.58 1315.20,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1290.00,1110.00 Q 1297.32,1113.03 1303.20,1110.00 Q 1297.32,1106.97 1290.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,1110.00 Q 1293.03,1117.32 1299.33,1119.33 Q 1297.32,1113.03 1290.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,1110.00 Q 1286.97,1117.32 1290.00,1123.20 Q 1293.03,1117.32 1290.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,1110.00 Q 1282.68,1113.03 1280.67,1119.33 Q 1286.97,1117.32 1290.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,1110.00 Q 1282.68,1106.97 1276.80,1110.00 Q 1282.68,1113.03 1290.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,1110.00 Q 1286.97,1102.68 1280.67,1100.67 Q 1282.68,1106.97 1290.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,1110.00 Q 1293.03,1102.68 1290.00,1096.80 Q 1286.97,1102.68 1290.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,1110.00 Q 1297.32,1106.97 1299.33,1100.67 Q 1293.03,1102.68 1290.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1290.00,1110.00 Q 1290.93,1113.48 1295.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,1110.00 Q 1286.52,1110.93 1284.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,1110.00 Q 1289.07,1106.52 1284.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1290.00,1110.00 Q 1293.48,1109.07 1295.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1290.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1274.88,1110.00 C 1281.28,1103.60 1288.14,1096.74 1290.00,1094.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1305.12,1110.00 C 1298.72,1116.40 1291.86,1123.26 1290.00,1125.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1350.00,1135.20 C 1339.02,1124.22 1328.22,1113.42 1324.80,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,1084.80 C 1360.98,1095.78 1371.78,1106.58 1375.20,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.8"><path d="M 1350.00,1110.00 Q 1357.32,1113.03 1363.20,1110.00 Q 1357.32,1106.97 1350.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,1110.00 Q 1353.03,1117.32 1359.33,1119.33 Q 1357.32,1113.03 1350.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,1110.00 Q 1346.97,1117.32 1350.00,1123.20 Q 1353.03,1117.32 1350.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,1110.00 Q 1342.68,1113.03 1340.67,1119.33 Q 1346.97,1117.32 1350.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,1110.00 Q 1342.68,1106.97 1336.80,1110.00 Q 1342.68,1113.03 1350.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,1110.00 Q 1346.97,1102.68 1340.67,1100.67 Q 1342.68,1106.97 1350.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,1110.00 Q 1353.03,1102.68 1350.00,1096.80 Q 1346.97,1102.68 1350.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,1110.00 Q 1357.32,1106.97 1359.33,1100.67 Q 1353.03,1102.68 1350.00,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.8999999999999999" /><path d="M 1350.00,1110.00 Q 1350.93,1113.48 1355.09,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,1110.00 Q 1346.52,1110.93 1344.91,1115.09" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,1110.00 Q 1349.07,1106.52 1344.91,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><path d="M 1350.00,1110.00 Q 1353.48,1109.07 1355.09,1104.91" fill="none" stroke="#000000" stroke-linecap="round" stroke-width="0.6" /><circle cx="1350.0" cy="1110.0" fill="none" opacity="0.6" r="4.8" stroke="#000000" stroke-width="0.72" /></g><g opacity="0.18"><path d="M 1334.88,1110.00 C 1341.28,1103.60 1348.14,1096.74 1350.00,1094.88" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1365.12,1110.00 C 1358.72,1116.40 1351.86,1123.26 1350.00,1125.12" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 175.20,1170.00 C 164.22,1180.98 153.42,1191.78 150.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 124.80,1170.00 C 135.78,1159.02 146.58,1148.22 150.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 150.00,1185.12 C 143.60,1178.72 136.74,1171.86 134.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,1154.88 C 156.40,1161.28 163.26,1168.14 165.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 184.80,1170.00 C 195.78,1159.02 206.58,1148.22 210.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 235.20,1170.00 C 224.22,1180.98 213.42,1191.78 210.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,1154.88 C 216.40,1161.28 223.26,1168.14 225.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,1185.12 C 203.60,1178.72 196.74,1171.86 194.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 244.80,1170.00 C 255.78,1159.02 266.58,1148.22 270.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 295.20,1170.00 C 284.22,1180.98 273.42,1191.78 270.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 270.00,1154.88 C 276.40,1161.28 283.26,1168.14 285.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,1185.12 C 263.60,1178.72 256.74,1171.86 254.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,1170.00 C 315.78,1159.02 326.58,1148.22 330.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,1170.00 C 344.22,1180.98 333.42,1191.78 330.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 330.00,1154.88 C 336.40,1161.28 343.26,1168.14 345.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,1185.12 C 323.60,1178.72 316.74,1171.86 314.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,1170.00 C 375.78,1159.02 386.58,1148.22 390.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,1170.00 C 404.22,1180.98 393.42,1191.78 390.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 390.00,1154.88 C 396.40,1161.28 403.26,1168.14 405.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,1185.12 C 383.60,1178.72 376.74,1171.86 374.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 424.80,1170.00 C 435.78,1159.02 446.58,1148.22 450.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 475.20,1170.00 C 464.22,1180.98 453.42,1191.78 450.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 450.00,1154.88 C 456.40,1161.28 463.26,1168.14 465.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,1185.12 C 443.60,1178.72 436.74,1171.86 434.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 484.80,1170.00 C 495.78,1159.02 506.58,1148.22 510.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 535.20,1170.00 C 524.22,1180.98 513.42,1191.78 510.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 510.00,1154.88 C 516.40,1161.28 523.26,1168.14 525.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,1185.12 C 503.60,1178.72 496.74,1171.86 494.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,1170.00 C 555.78,1159.02 566.58,1148.22 570.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,1170.00 C 584.22,1180.98 573.42,1191.78 570.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 570.00,1154.88 C 576.40,1161.28 583.26,1168.14 585.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,1185.12 C 563.60,1178.72 556.74,1171.86 554.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,1170.00 C 615.78,1159.02 626.58,1148.22 630.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,1170.00 C 644.22,1180.98 633.42,1191.78 630.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,1154.88 C 636.40,1161.28 643.26,1168.14 645.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,1185.12 C 623.60,1178.72 616.74,1171.86 614.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 664.80,1170.00 C 675.78,1159.02 686.58,1148.22 690.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 715.20,1170.00 C 704.22,1180.98 693.42,1191.78 690.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 690.00,1154.88 C 696.40,1161.28 703.26,1168.14 705.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,1185.12 C 683.60,1178.72 676.74,1171.86 674.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 724.80,1170.00 C 735.78,1159.02 746.58,1148.22 750.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 775.20,1170.00 C 764.22,1180.98 753.42,1191.78 750.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,1154.88 C 756.40,1161.28 763.26,1168.14 765.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,1185.12 C 743.60,1178.72 736.74,1171.86 734.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 784.80,1170.00 C 795.78,1159.02 806.58,1148.22 810.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 835.20,1170.00 C 824.22,1180.98 813.42,1191.78 810.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,1154.88 C 816.40,1161.28 823.26,1168.14 825.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,1185.12 C 803.60,1178.72 796.74,1171.86 794.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 844.80,1170.00 C 855.78,1159.02 866.58,1148.22 870.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 895.20,1170.00 C 884.22,1180.98 873.42,1191.78 870.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 870.00,1154.88 C 876.40,1161.28 883.26,1168.14 885.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,1185.12 C 863.60,1178.72 856.74,1171.86 854.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 904.80,1170.00 C 915.78,1159.02 926.58,1148.22 930.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 955.20,1170.00 C 944.22,1180.98 933.42,1191.78 930.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 930.00,1154.88 C 936.40,1161.28 943.26,1168.14 945.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,1185.12 C 923.60,1178.72 916.74,1171.86 914.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 964.80,1170.00 C 975.78,1159.02 986.58,1148.22 990.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1015.20,1170.00 C 1004.22,1180.98 993.42,1191.78 990.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 990.00,1154.88 C 996.40,1161.28 1003.26,1168.14 1005.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,1185.12 C 983.60,1178.72 976.74,1171.86 974.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,1170.00 C 1035.78,1159.02 1046.58,1148.22 1050.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,1170.00 C 1064.22,1180.98 1053.42,1191.78 1050.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,1154.88 C 1056.40,1161.28 1063.26,1168.14 1065.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,1185.12 C 1043.60,1178.72 1036.74,1171.86 1034.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1084.80,1170.00 C 1095.78,1159.02 1106.58,1148.22 1110.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1135.20,1170.00 C 1124.22,1180.98 1113.42,1191.78 1110.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1110.00,1154.88 C 1116.40,1161.28 1123.26,1168.14 1125.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,1185.12 C 1103.60,1178.72 1096.74,1171.86 1094.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1144.80,1170.00 C 1155.78,1159.02 1166.58,1148.22 1170.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1195.20,1170.00 C 1184.22,1180.98 1173.42,1191.78 1170.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1170.00,1154.88 C 1176.40,1161.28 1183.26,1168.14 1185.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,1185.12 C 1163.60,1178.72 1156.74,1171.86 1154.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1204.80,1170.00 C 1215.78,1159.02 1226.58,1148.22 1230.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1255.20,1170.00 C 1244.22,1180.98 1233.42,1191.78 1230.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1230.00,1154.88 C 1236.40,1161.28 1243.26,1168.14 1245.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,1185.12 C 1223.60,1178.72 1216.74,1171.86 1214.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1264.80,1170.00 C 1275.78,1159.02 1286.58,1148.22 1290.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1315.20,1170.00 C 1304.22,1180.98 1293.42,1191.78 1290.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1290.00,1154.88 C 1296.40,1161.28 1303.26,1168.14 1305.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,1185.12 C 1283.60,1178.72 1276.74,1171.86 1274.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1324.80,1170.00 C 1335.78,1159.02 1346.58,1148.22 1350.00,1144.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1375.20,1170.00 C 1364.22,1180.98 1353.42,1191.78 1350.00,1195.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,1154.88 C 1356.40,1161.28 1363.26,1168.14 1365.12,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,1185.12 C 1343.60,1178.72 1336.74,1171.86 1334.88,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 124.80,1230.00 C 135.78,1219.02 146.58,1208.22 150.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 175.20,1230.00 C 164.22,1240.98 153.42,1251.78 150.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 150.00,1214.88 C 156.40,1221.28 163.26,1228.14 165.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,1245.12 C 143.60,1238.72 136.74,1231.86 134.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 184.80,1230.00 C 195.78,1219.02 206.58,1208.22 210.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 235.20,1230.00 C 224.22,1240.98 213.42,1251.78 210.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,1214.88 C 216.40,1221.28 223.26,1228.14 225.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,1245.12 C 203.60,1238.72 196.74,1231.86 194.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 244.80,1230.00 C 255.78,1219.02 266.58,1208.22 270.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 295.20,1230.00 C 284.22,1240.98 273.42,1251.78 270.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 270.00,1214.88 C 276.40,1221.28 283.26,1228.14 285.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,1245.12 C 263.60,1238.72 256.74,1231.86 254.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,1230.00 C 315.78,1219.02 326.58,1208.22 330.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,1230.00 C 344.22,1240.98 333.42,1251.78 330.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 330.00,1214.88 C 336.40,1221.28 343.26,1228.14 345.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,1245.12 C 323.60,1238.72 316.74,1231.86 314.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,1230.00 C 375.78,1219.02 386.58,1208.22 390.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,1230.00 C 404.22,1240.98 393.42,1251.78 390.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 390.00,1214.88 C 396.40,1221.28 403.26,1228.14 405.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,1245.12 C 383.60,1238.72 376.74,1231.86 374.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 424.80,1230.00 C 435.78,1219.02 446.58,1208.22 450.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 475.20,1230.00 C 464.22,1240.98 453.42,1251.78 450.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 450.00,1214.88 C 456.40,1221.28 463.26,1228.14 465.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,1245.12 C 443.60,1238.72 436.74,1231.86 434.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 484.80,1230.00 C 495.78,1219.02 506.58,1208.22 510.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 535.20,1230.00 C 524.22,1240.98 513.42,1251.78 510.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 510.00,1214.88 C 516.40,1221.28 523.26,1228.14 525.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,1245.12 C 503.60,1238.72 496.74,1231.86 494.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,1230.00 C 555.78,1219.02 566.58,1208.22 570.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,1230.00 C 584.22,1240.98 573.42,1251.78 570.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 570.00,1214.88 C 576.40,1221.28 583.26,1228.14 585.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,1245.12 C 563.60,1238.72 556.74,1231.86 554.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,1230.00 C 615.78,1219.02 626.58,1208.22 630.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,1230.00 C 644.22,1240.98 633.42,1251.78 630.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,1214.88 C 636.40,1221.28 643.26,1228.14 645.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,1245.12 C 623.60,1238.72 616.74,1231.86 614.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 664.80,1230.00 C 675.78,1219.02 686.58,1208.22 690.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 715.20,1230.00 C 704.22,1240.98 693.42,1251.78 690.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 690.00,1214.88 C 696.40,1221.28 703.26,1228.14 705.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,1245.12 C 683.60,1238.72 676.74,1231.86 674.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 724.80,1230.00 C 735.78,1219.02 746.58,1208.22 750.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 775.20,1230.00 C 764.22,1240.98 753.42,1251.78 750.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,1214.88 C 756.40,1221.28 763.26,1228.14 765.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,1245.12 C 743.60,1238.72 736.74,1231.86 734.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 784.80,1230.00 C 795.78,1219.02 806.58,1208.22 810.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 835.20,1230.00 C 824.22,1240.98 813.42,1251.78 810.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,1214.88 C 816.40,1221.28 823.26,1228.14 825.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,1245.12 C 803.60,1238.72 796.74,1231.86 794.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 844.80,1230.00 C 855.78,1219.02 866.58,1208.22 870.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 895.20,1230.00 C 884.22,1240.98 873.42,1251.78 870.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 870.00,1214.88 C 876.40,1221.28 883.26,1228.14 885.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,1245.12 C 863.60,1238.72 856.74,1231.86 854.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 904.80,1230.00 C 915.78,1219.02 926.58,1208.22 930.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 955.20,1230.00 C 944.22,1240.98 933.42,1251.78 930.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 930.00,1214.88 C 936.40,1221.28 943.26,1228.14 945.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,1245.12 C 923.60,1238.72 916.74,1231.86 914.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 964.80,1230.00 C 975.78,1219.02 986.58,1208.22 990.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1015.20,1230.00 C 1004.22,1240.98 993.42,1251.78 990.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 990.00,1214.88 C 996.40,1221.28 1003.26,1228.14 1005.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,1245.12 C 983.60,1238.72 976.74,1231.86 974.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,1230.00 C 1035.78,1219.02 1046.58,1208.22 1050.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,1230.00 C 1064.22,1240.98 1053.42,1251.78 1050.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,1214.88 C 1056.40,1221.28 1063.26,1228.14 1065.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,1245.12 C 1043.60,1238.72 1036.74,1231.86 1034.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1084.80,1230.00 C 1095.78,1219.02 1106.58,1208.22 1110.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1135.20,1230.00 C 1124.22,1240.98 1113.42,1251.78 1110.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1110.00,1214.88 C 1116.40,1221.28 1123.26,1228.14 1125.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,1245.12 C 1103.60,1238.72 1096.74,1231.86 1094.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1144.80,1230.00 C 1155.78,1219.02 1166.58,1208.22 1170.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1195.20,1230.00 C 1184.22,1240.98 1173.42,1251.78 1170.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1170.00,1214.88 C 1176.40,1221.28 1183.26,1228.14 1185.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,1245.12 C 1163.60,1238.72 1156.74,1231.86 1154.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1204.80,1230.00 C 1215.78,1219.02 1226.58,1208.22 1230.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1255.20,1230.00 C 1244.22,1240.98 1233.42,1251.78 1230.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1230.00,1214.88 C 1236.40,1221.28 1243.26,1228.14 1245.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,1245.12 C 1223.60,1238.72 1216.74,1231.86 1214.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1264.80,1230.00 C 1275.78,1219.02 1286.58,1208.22 1290.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1315.20,1230.00 C 1304.22,1240.98 1293.42,1251.78 1290.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1290.00,1214.88 C 1296.40,1221.28 1303.26,1228.14 1305.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,1245.12 C 1283.60,1238.72 1276.74,1231.86 1274.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1324.80,1230.00 C 1335.78,1219.02 1346.58,1208.22 1350.00,1204.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1375.20,1230.00 C 1364.22,1240.98 1353.42,1251.78 1350.00,1255.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,1214.88 C 1356.40,1221.28 1363.26,1228.14 1365.12,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,1245.12 C 1343.60,1238.72 1336.74,1231.86 1334.88,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 124.80,1290.00 C 135.78,1279.02 146.58,1268.22 150.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 175.20,1290.00 C 164.22,1300.98 153.42,1311.78 150.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 150.00,1274.88 C 156.40,1281.28 163.26,1288.14 165.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,1305.12 C 143.60,1298.72 136.74,1291.86 134.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 184.80,1290.00 C 195.78,1279.02 206.58,1268.22 210.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 235.20,1290.00 C 224.22,1300.98 213.42,1311.78 210.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,1274.88 C 216.40,1281.28 223.26,1288.14 225.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,1305.12 C 203.60,1298.72 196.74,1291.86 194.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 244.80,1290.00 C 255.78,1279.02 266.58,1268.22 270.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 295.20,1290.00 C 284.22,1300.98 273.42,1311.78 270.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 270.00,1274.88 C 276.40,1281.28 283.26,1288.14 285.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,1305.12 C 263.60,1298.72 256.74,1291.86 254.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,1290.00 C 315.78,1279.02 326.58,1268.22 330.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,1290.00 C 344.22,1300.98 333.42,1311.78 330.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 330.00,1274.88 C 336.40,1281.28 343.26,1288.14 345.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,1305.12 C 323.60,1298.72 316.74,1291.86 314.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,1290.00 C 375.78,1279.02 386.58,1268.22 390.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,1290.00 C 404.22,1300.98 393.42,1311.78 390.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 390.00,1274.88 C 396.40,1281.28 403.26,1288.14 405.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,1305.12 C 383.60,1298.72 376.74,1291.86 374.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 424.80,1290.00 C 435.78,1279.02 446.58,1268.22 450.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 475.20,1290.00 C 464.22,1300.98 453.42,1311.78 450.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 450.00,1274.88 C 456.40,1281.28 463.26,1288.14 465.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,1305.12 C 443.60,1298.72 436.74,1291.86 434.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 484.80,1290.00 C 495.78,1279.02 506.58,1268.22 510.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 535.20,1290.00 C 524.22,1300.98 513.42,1311.78 510.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 510.00,1274.88 C 516.40,1281.28 523.26,1288.14 525.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,1305.12 C 503.60,1298.72 496.74,1291.86 494.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,1290.00 C 555.78,1279.02 566.58,1268.22 570.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,1290.00 C 584.22,1300.98 573.42,1311.78 570.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 570.00,1274.88 C 576.40,1281.28 583.26,1288.14 585.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,1305.12 C 563.60,1298.72 556.74,1291.86 554.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,1290.00 C 615.78,1279.02 626.58,1268.22 630.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,1290.00 C 644.22,1300.98 633.42,1311.78 630.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,1274.88 C 636.40,1281.28 643.26,1288.14 645.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,1305.12 C 623.60,1298.72 616.74,1291.86 614.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 664.80,1290.00 C 675.78,1279.02 686.58,1268.22 690.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 715.20,1290.00 C 704.22,1300.98 693.42,1311.78 690.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 690.00,1274.88 C 696.40,1281.28 703.26,1288.14 705.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,1305.12 C 683.60,1298.72 676.74,1291.86 674.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 724.80,1290.00 C 735.78,1279.02 746.58,1268.22 750.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 775.20,1290.00 C 764.22,1300.98 753.42,1311.78 750.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,1274.88 C 756.40,1281.28 763.26,1288.14 765.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,1305.12 C 743.60,1298.72 736.74,1291.86 734.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 784.80,1290.00 C 795.78,1279.02 806.58,1268.22 810.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 835.20,1290.00 C 824.22,1300.98 813.42,1311.78 810.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,1274.88 C 816.40,1281.28 823.26,1288.14 825.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,1305.12 C 803.60,1298.72 796.74,1291.86 794.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 844.80,1290.00 C 855.78,1279.02 866.58,1268.22 870.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 895.20,1290.00 C 884.22,1300.98 873.42,1311.78 870.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 870.00,1274.88 C 876.40,1281.28 883.26,1288.14 885.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,1305.12 C 863.60,1298.72 856.74,1291.86 854.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 904.80,1290.00 C 915.78,1279.02 926.58,1268.22 930.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 955.20,1290.00 C 944.22,1300.98 933.42,1311.78 930.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 930.00,1274.88 C 936.40,1281.28 943.26,1288.14 945.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,1305.12 C 923.60,1298.72 916.74,1291.86 914.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 964.80,1290.00 C 975.78,1279.02 986.58,1268.22 990.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1015.20,1290.00 C 1004.22,1300.98 993.42,1311.78 990.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 990.00,1274.88 C 996.40,1281.28 1003.26,1288.14 1005.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,1305.12 C 983.60,1298.72 976.74,1291.86 974.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,1290.00 C 1035.78,1279.02 1046.58,1268.22 1050.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,1290.00 C 1064.22,1300.98 1053.42,1311.78 1050.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,1274.88 C 1056.40,1281.28 1063.26,1288.14 1065.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,1305.12 C 1043.60,1298.72 1036.74,1291.86 1034.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1084.80,1290.00 C 1095.78,1279.02 1106.58,1268.22 1110.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1135.20,1290.00 C 1124.22,1300.98 1113.42,1311.78 1110.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1110.00,1274.88 C 1116.40,1281.28 1123.26,1288.14 1125.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,1305.12 C 1103.60,1298.72 1096.74,1291.86 1094.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1144.80,1290.00 C 1155.78,1279.02 1166.58,1268.22 1170.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1195.20,1290.00 C 1184.22,1300.98 1173.42,1311.78 1170.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1170.00,1274.88 C 1176.40,1281.28 1183.26,1288.14 1185.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,1305.12 C 1163.60,1298.72 1156.74,1291.86 1154.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1204.80,1290.00 C 1215.78,1279.02 1226.58,1268.22 1230.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1255.20,1290.00 C 1244.22,1300.98 1233.42,1311.78 1230.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1230.00,1274.88 C 1236.40,1281.28 1243.26,1288.14 1245.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,1305.12 C 1223.60,1298.72 1216.74,1291.86 1214.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1264.80,1290.00 C 1275.78,1279.02 1286.58,1268.22 1290.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1315.20,1290.00 C 1304.22,1300.98 1293.42,1311.78 1290.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1290.00,1274.88 C 1296.40,1281.28 1303.26,1288.14 1305.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,1305.12 C 1283.60,1298.72 1276.74,1291.86 1274.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1324.80,1290.00 C 1335.78,1279.02 1346.58,1268.22 1350.00,1264.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1375.20,1290.00 C 1364.22,1300.98 1353.42,1311.78 1350.00,1315.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,1274.88 C 1356.40,1281.28 1363.26,1288.14 1365.12,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,1305.12 C 1343.60,1298.72 1336.74,1291.86 1334.88,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 124.80,1350.00 C 135.78,1339.02 146.58,1328.22 150.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 175.20,1350.00 C 164.22,1360.98 153.42,1371.78 150.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 150.00,1334.88 C 156.40,1341.28 163.26,1348.14 165.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 150.00,1365.12 C 143.60,1358.72 136.74,1351.86 134.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 184.80,1350.00 C 195.78,1339.02 206.58,1328.22 210.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 235.20,1350.00 C 224.22,1360.98 213.42,1371.78 210.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 210.00,1334.88 C 216.40,1341.28 223.26,1348.14 225.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 210.00,1365.12 C 203.60,1358.72 196.74,1351.86 194.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 244.80,1350.00 C 255.78,1339.02 266.58,1328.22 270.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 295.20,1350.00 C 284.22,1360.98 273.42,1371.78 270.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 270.00,1334.88 C 276.40,1341.28 283.26,1348.14 285.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 270.00,1365.12 C 263.60,1358.72 256.74,1351.86 254.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 304.80,1350.00 C 315.78,1339.02 326.58,1328.22 330.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 355.20,1350.00 C 344.22,1360.98 333.42,1371.78 330.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 330.00,1334.88 C 336.40,1341.28 343.26,1348.14 345.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 330.00,1365.12 C 323.60,1358.72 316.74,1351.86 314.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 364.80,1350.00 C 375.78,1339.02 386.58,1328.22 390.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 415.20,1350.00 C 404.22,1360.98 393.42,1371.78 390.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 390.00,1334.88 C 396.40,1341.28 403.26,1348.14 405.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 390.00,1365.12 C 383.60,1358.72 376.74,1351.86 374.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 424.80,1350.00 C 435.78,1339.02 446.58,1328.22 450.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 475.20,1350.00 C 464.22,1360.98 453.42,1371.78 450.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 450.00,1334.88 C 456.40,1341.28 463.26,1348.14 465.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 450.00,1365.12 C 443.60,1358.72 436.74,1351.86 434.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 484.80,1350.00 C 495.78,1339.02 506.58,1328.22 510.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 535.20,1350.00 C 524.22,1360.98 513.42,1371.78 510.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 510.00,1334.88 C 516.40,1341.28 523.26,1348.14 525.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 510.00,1365.12 C 503.60,1358.72 496.74,1351.86 494.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 544.80,1350.00 C 555.78,1339.02 566.58,1328.22 570.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 595.20,1350.00 C 584.22,1360.98 573.42,1371.78 570.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 570.00,1334.88 C 576.40,1341.28 583.26,1348.14 585.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 570.00,1365.12 C 563.60,1358.72 556.74,1351.86 554.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 604.80,1350.00 C 615.78,1339.02 626.58,1328.22 630.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 655.20,1350.00 C 644.22,1360.98 633.42,1371.78 630.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 630.00,1334.88 C 636.40,1341.28 643.26,1348.14 645.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 630.00,1365.12 C 623.60,1358.72 616.74,1351.86 614.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 664.80,1350.00 C 675.78,1339.02 686.58,1328.22 690.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 715.20,1350.00 C 704.22,1360.98 693.42,1371.78 690.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 690.00,1334.88 C 696.40,1341.28 703.26,1348.14 705.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 690.00,1365.12 C 683.60,1358.72 676.74,1351.86 674.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 724.80,1350.00 C 735.78,1339.02 746.58,1328.22 750.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 775.20,1350.00 C 764.22,1360.98 753.42,1371.78 750.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 750.00,1334.88 C 756.40,1341.28 763.26,1348.14 765.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 750.00,1365.12 C 743.60,1358.72 736.74,1351.86 734.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 784.80,1350.00 C 795.78,1339.02 806.58,1328.22 810.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 835.20,1350.00 C 824.22,1360.98 813.42,1371.78 810.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 810.00,1334.88 C 816.40,1341.28 823.26,1348.14 825.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 810.00,1365.12 C 803.60,1358.72 796.74,1351.86 794.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 844.80,1350.00 C 855.78,1339.02 866.58,1328.22 870.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 895.20,1350.00 C 884.22,1360.98 873.42,1371.78 870.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 870.00,1334.88 C 876.40,1341.28 883.26,1348.14 885.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 870.00,1365.12 C 863.60,1358.72 856.74,1351.86 854.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 904.80,1350.00 C 915.78,1339.02 926.58,1328.22 930.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 955.20,1350.00 C 944.22,1360.98 933.42,1371.78 930.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 930.00,1334.88 C 936.40,1341.28 943.26,1348.14 945.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 930.00,1365.12 C 923.60,1358.72 916.74,1351.86 914.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 964.80,1350.00 C 975.78,1339.02 986.58,1328.22 990.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1015.20,1350.00 C 1004.22,1360.98 993.42,1371.78 990.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 990.00,1334.88 C 996.40,1341.28 1003.26,1348.14 1005.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 990.00,1365.12 C 983.60,1358.72 976.74,1351.86 974.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1024.80,1350.00 C 1035.78,1339.02 1046.58,1328.22 1050.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1075.20,1350.00 C 1064.22,1360.98 1053.42,1371.78 1050.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1050.00,1334.88 C 1056.40,1341.28 1063.26,1348.14 1065.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1050.00,1365.12 C 1043.60,1358.72 1036.74,1351.86 1034.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1084.80,1350.00 C 1095.78,1339.02 1106.58,1328.22 1110.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1135.20,1350.00 C 1124.22,1360.98 1113.42,1371.78 1110.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1110.00,1334.88 C 1116.40,1341.28 1123.26,1348.14 1125.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1110.00,1365.12 C 1103.60,1358.72 1096.74,1351.86 1094.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1144.80,1350.00 C 1155.78,1339.02 1166.58,1328.22 1170.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1195.20,1350.00 C 1184.22,1360.98 1173.42,1371.78 1170.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1170.00,1334.88 C 1176.40,1341.28 1183.26,1348.14 1185.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1170.00,1365.12 C 1163.60,1358.72 1156.74,1351.86 1154.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1204.80,1350.00 C 1215.78,1339.02 1226.58,1328.22 1230.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1255.20,1350.00 C 1244.22,1360.98 1233.42,1371.78 1230.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1230.00,1334.88 C 1236.40,1341.28 1243.26,1348.14 1245.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1230.00,1365.12 C 1223.60,1358.72 1216.74,1351.86 1214.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1264.80,1350.00 C 1275.78,1339.02 1286.58,1328.22 1290.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1315.20,1350.00 C 1304.22,1360.98 1293.42,1371.78 1290.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1290.00,1334.88 C 1296.40,1341.28 1303.26,1348.14 1305.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1290.00,1365.12 C 1283.60,1358.72 1276.74,1351.86 1274.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 1324.80,1350.00 C 1335.78,1339.02 1346.58,1328.22 1350.00,1324.80" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1375.20,1350.00 C 1364.22,1360.98 1353.42,1371.78 1350.00,1375.20" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><g opacity="0.18"><path d="M 1350.00,1334.88 C 1356.40,1341.28 1363.26,1348.14 1365.12,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /><path d="M 1350.00,1365.12 C 1343.60,1358.72 1336.74,1351.86 1334.88,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.0" /></g><path d="M 164.70,150.00 C 171.00,161.76 179.40,161.76 185.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,150.00 C 171.00,161.76 179.40,161.76 185.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,150.00 C 171.00,161.76 179.40,161.76 185.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,150.00 C 231.00,161.76 239.40,161.76 245.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,150.00 C 231.00,161.76 239.40,161.76 245.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,150.00 C 231.00,161.76 239.40,161.76 245.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,150.00 C 291.00,161.76 299.40,161.76 305.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,150.00 C 291.00,161.76 299.40,161.76 305.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,150.00 C 291.00,161.76 299.40,161.76 305.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,150.00 C 351.00,161.76 359.40,161.76 365.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,150.00 C 351.00,161.76 359.40,161.76 365.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,150.00 C 351.00,161.76 359.40,161.76 365.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,150.00 C 411.00,161.76 419.40,161.76 425.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,150.00 C 411.00,161.76 419.40,161.76 425.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,150.00 C 411.00,161.76 419.40,161.76 425.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,150.00 C 471.00,161.76 479.40,161.76 485.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,150.00 C 471.00,161.76 479.40,161.76 485.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,150.00 C 471.00,161.76 479.40,161.76 485.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,150.00 C 531.00,161.76 539.40,161.76 545.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,150.00 C 531.00,161.76 539.40,161.76 545.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,150.00 C 531.00,161.76 539.40,161.76 545.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,150.00 C 591.00,161.76 599.40,161.76 605.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,150.00 C 591.00,161.76 599.40,161.76 605.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,150.00 C 591.00,161.76 599.40,161.76 605.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,150.00 C 651.00,161.76 659.40,161.76 665.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,150.00 C 651.00,161.76 659.40,161.76 665.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,150.00 C 651.00,161.76 659.40,161.76 665.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,150.00 C 711.00,161.76 719.40,161.76 725.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,150.00 C 711.00,161.76 719.40,161.76 725.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,150.00 C 711.00,161.76 719.40,161.76 725.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,150.00 C 771.00,161.76 779.40,161.76 785.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,150.00 C 771.00,161.76 779.40,161.76 785.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,150.00 C 771.00,161.76 779.40,161.76 785.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,150.00 C 831.00,161.76 839.40,161.76 845.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,150.00 C 831.00,161.76 839.40,161.76 845.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,150.00 C 831.00,161.76 839.40,161.76 845.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,150.00 C 891.00,161.76 899.40,161.76 905.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,150.00 C 891.00,161.76 899.40,161.76 905.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,150.00 C 891.00,161.76 899.40,161.76 905.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,150.00 C 951.00,161.76 959.40,161.76 965.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,150.00 C 951.00,161.76 959.40,161.76 965.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,150.00 C 951.00,161.76 959.40,161.76 965.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,150.00 C 1011.00,161.76 1019.40,161.76 1025.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,150.00 C 1011.00,161.76 1019.40,161.76 1025.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,150.00 C 1011.00,161.76 1019.40,161.76 1025.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,150.00 C 1071.00,161.76 1079.40,161.76 1085.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,150.00 C 1071.00,161.76 1079.40,161.76 1085.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,150.00 C 1071.00,161.76 1079.40,161.76 1085.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,150.00 C 1131.00,161.76 1139.40,161.76 1145.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,150.00 C 1131.00,161.76 1139.40,161.76 1145.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,150.00 C 1131.00,161.76 1139.40,161.76 1145.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,150.00 C 1191.00,161.76 1199.40,161.76 1205.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,150.00 C 1191.00,161.76 1199.40,161.76 1205.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,150.00 C 1191.00,161.76 1199.40,161.76 1205.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,150.00 C 1251.00,161.76 1259.40,161.76 1265.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,150.00 C 1251.00,161.76 1259.40,161.76 1265.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,150.00 C 1251.00,161.76 1259.40,161.76 1265.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,150.00 C 1311.00,161.76 1319.40,161.76 1325.70,150.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,150.00 C 1311.00,161.76 1319.40,161.76 1325.70,150.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,150.00 C 1311.00,161.76 1319.40,161.76 1325.70,150.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,210.00 C 171.00,221.76 179.40,221.76 185.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,210.00 C 171.00,221.76 179.40,221.76 185.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,210.00 C 171.00,221.76 179.40,221.76 185.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,210.00 C 231.00,221.76 239.40,221.76 245.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,210.00 C 231.00,221.76 239.40,221.76 245.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,210.00 C 231.00,221.76 239.40,221.76 245.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,210.00 C 291.00,221.76 299.40,221.76 305.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,210.00 C 291.00,221.76 299.40,221.76 305.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,210.00 C 291.00,221.76 299.40,221.76 305.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,210.00 C 351.00,221.76 359.40,221.76 365.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,210.00 C 351.00,221.76 359.40,221.76 365.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,210.00 C 351.00,221.76 359.40,221.76 365.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,210.00 C 411.00,221.76 419.40,221.76 425.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,210.00 C 411.00,221.76 419.40,221.76 425.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,210.00 C 411.00,221.76 419.40,221.76 425.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,210.00 C 471.00,221.76 479.40,221.76 485.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,210.00 C 471.00,221.76 479.40,221.76 485.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,210.00 C 471.00,221.76 479.40,221.76 485.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,210.00 C 531.00,221.76 539.40,221.76 545.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,210.00 C 531.00,221.76 539.40,221.76 545.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,210.00 C 531.00,221.76 539.40,221.76 545.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,210.00 C 591.00,221.76 599.40,221.76 605.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,210.00 C 591.00,221.76 599.40,221.76 605.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,210.00 C 591.00,221.76 599.40,221.76 605.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,210.00 C 651.00,221.76 659.40,221.76 665.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,210.00 C 651.00,221.76 659.40,221.76 665.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,210.00 C 651.00,221.76 659.40,221.76 665.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,210.00 C 711.00,221.76 719.40,221.76 725.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,210.00 C 711.00,221.76 719.40,221.76 725.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,210.00 C 711.00,221.76 719.40,221.76 725.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,210.00 C 771.00,221.76 779.40,221.76 785.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,210.00 C 771.00,221.76 779.40,221.76 785.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,210.00 C 771.00,221.76 779.40,221.76 785.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,210.00 C 831.00,221.76 839.40,221.76 845.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,210.00 C 831.00,221.76 839.40,221.76 845.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,210.00 C 831.00,221.76 839.40,221.76 845.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,210.00 C 891.00,221.76 899.40,221.76 905.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,210.00 C 891.00,221.76 899.40,221.76 905.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,210.00 C 891.00,221.76 899.40,221.76 905.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,210.00 C 951.00,221.76 959.40,221.76 965.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,210.00 C 951.00,221.76 959.40,221.76 965.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,210.00 C 951.00,221.76 959.40,221.76 965.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,210.00 C 1011.00,221.76 1019.40,221.76 1025.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,210.00 C 1011.00,221.76 1019.40,221.76 1025.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,210.00 C 1011.00,221.76 1019.40,221.76 1025.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,210.00 C 1071.00,221.76 1079.40,221.76 1085.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,210.00 C 1071.00,221.76 1079.40,221.76 1085.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,210.00 C 1071.00,221.76 1079.40,221.76 1085.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,210.00 C 1131.00,221.76 1139.40,221.76 1145.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,210.00 C 1131.00,221.76 1139.40,221.76 1145.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,210.00 C 1131.00,221.76 1139.40,221.76 1145.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,210.00 C 1191.00,221.76 1199.40,221.76 1205.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,210.00 C 1191.00,221.76 1199.40,221.76 1205.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,210.00 C 1191.00,221.76 1199.40,221.76 1205.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,210.00 C 1251.00,221.76 1259.40,221.76 1265.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,210.00 C 1251.00,221.76 1259.40,221.76 1265.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,210.00 C 1251.00,221.76 1259.40,221.76 1265.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,210.00 C 1311.00,221.76 1319.40,221.76 1325.70,210.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,210.00 C 1311.00,221.76 1319.40,221.76 1325.70,210.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,210.00 C 1311.00,221.76 1319.40,221.76 1325.70,210.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,270.00 C 171.00,281.76 179.40,281.76 185.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,270.00 C 171.00,281.76 179.40,281.76 185.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,270.00 C 171.00,281.76 179.40,281.76 185.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,270.00 C 231.00,281.76 239.40,281.76 245.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,270.00 C 231.00,281.76 239.40,281.76 245.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,270.00 C 231.00,281.76 239.40,281.76 245.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,270.00 C 291.00,281.76 299.40,281.76 305.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,270.00 C 291.00,281.76 299.40,281.76 305.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,270.00 C 291.00,281.76 299.40,281.76 305.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,270.00 C 351.00,281.76 359.40,281.76 365.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,270.00 C 351.00,281.76 359.40,281.76 365.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,270.00 C 351.00,281.76 359.40,281.76 365.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,270.00 C 411.00,281.76 419.40,281.76 425.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,270.00 C 411.00,281.76 419.40,281.76 425.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,270.00 C 411.00,281.76 419.40,281.76 425.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,270.00 C 471.00,281.76 479.40,281.76 485.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,270.00 C 471.00,281.76 479.40,281.76 485.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,270.00 C 471.00,281.76 479.40,281.76 485.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,270.00 C 531.00,281.76 539.40,281.76 545.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,270.00 C 531.00,281.76 539.40,281.76 545.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,270.00 C 531.00,281.76 539.40,281.76 545.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,270.00 C 591.00,281.76 599.40,281.76 605.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,270.00 C 591.00,281.76 599.40,281.76 605.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,270.00 C 591.00,281.76 599.40,281.76 605.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,270.00 C 651.00,281.76 659.40,281.76 665.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,270.00 C 651.00,281.76 659.40,281.76 665.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,270.00 C 651.00,281.76 659.40,281.76 665.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,270.00 C 711.00,281.76 719.40,281.76 725.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,270.00 C 711.00,281.76 719.40,281.76 725.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,270.00 C 711.00,281.76 719.40,281.76 725.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,270.00 C 771.00,281.76 779.40,281.76 785.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,270.00 C 771.00,281.76 779.40,281.76 785.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,270.00 C 771.00,281.76 779.40,281.76 785.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,270.00 C 831.00,281.76 839.40,281.76 845.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,270.00 C 831.00,281.76 839.40,281.76 845.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,270.00 C 831.00,281.76 839.40,281.76 845.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,270.00 C 891.00,281.76 899.40,281.76 905.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,270.00 C 891.00,281.76 899.40,281.76 905.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,270.00 C 891.00,281.76 899.40,281.76 905.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,270.00 C 951.00,281.76 959.40,281.76 965.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,270.00 C 951.00,281.76 959.40,281.76 965.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,270.00 C 951.00,281.76 959.40,281.76 965.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,270.00 C 1011.00,281.76 1019.40,281.76 1025.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,270.00 C 1011.00,281.76 1019.40,281.76 1025.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,270.00 C 1011.00,281.76 1019.40,281.76 1025.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,270.00 C 1071.00,281.76 1079.40,281.76 1085.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,270.00 C 1071.00,281.76 1079.40,281.76 1085.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,270.00 C 1071.00,281.76 1079.40,281.76 1085.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,270.00 C 1131.00,281.76 1139.40,281.76 1145.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,270.00 C 1131.00,281.76 1139.40,281.76 1145.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,270.00 C 1131.00,281.76 1139.40,281.76 1145.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,270.00 C 1191.00,281.76 1199.40,281.76 1205.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,270.00 C 1191.00,281.76 1199.40,281.76 1205.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,270.00 C 1191.00,281.76 1199.40,281.76 1205.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,270.00 C 1251.00,281.76 1259.40,281.76 1265.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,270.00 C 1251.00,281.76 1259.40,281.76 1265.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,270.00 C 1251.00,281.76 1259.40,281.76 1265.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,270.00 C 1311.00,281.76 1319.40,281.76 1325.70,270.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,270.00 C 1311.00,281.76 1319.40,281.76 1325.70,270.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,270.00 C 1311.00,281.76 1319.40,281.76 1325.70,270.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,330.00 C 171.00,341.76 179.40,341.76 185.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,330.00 C 171.00,341.76 179.40,341.76 185.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,330.00 C 171.00,341.76 179.40,341.76 185.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,330.00 C 231.00,341.76 239.40,341.76 245.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,330.00 C 231.00,341.76 239.40,341.76 245.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,330.00 C 231.00,341.76 239.40,341.76 245.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,330.00 C 291.00,341.76 299.40,341.76 305.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,330.00 C 291.00,341.76 299.40,341.76 305.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,330.00 C 291.00,341.76 299.40,341.76 305.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,330.00 C 351.00,341.76 359.40,341.76 365.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,330.00 C 351.00,341.76 359.40,341.76 365.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,330.00 C 351.00,341.76 359.40,341.76 365.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,330.00 C 411.00,341.76 419.40,341.76 425.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,330.00 C 411.00,341.76 419.40,341.76 425.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,330.00 C 411.00,341.76 419.40,341.76 425.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,330.00 C 471.00,341.76 479.40,341.76 485.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,330.00 C 471.00,341.76 479.40,341.76 485.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,330.00 C 471.00,341.76 479.40,341.76 485.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,330.00 C 531.00,341.76 539.40,341.76 545.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,330.00 C 531.00,341.76 539.40,341.76 545.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,330.00 C 531.00,341.76 539.40,341.76 545.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,330.00 C 591.00,341.76 599.40,341.76 605.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,330.00 C 591.00,341.76 599.40,341.76 605.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,330.00 C 591.00,341.76 599.40,341.76 605.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,330.00 C 651.00,341.76 659.40,341.76 665.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,330.00 C 651.00,341.76 659.40,341.76 665.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,330.00 C 651.00,341.76 659.40,341.76 665.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,330.00 C 711.00,341.76 719.40,341.76 725.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,330.00 C 711.00,341.76 719.40,341.76 725.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,330.00 C 711.00,341.76 719.40,341.76 725.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,330.00 C 771.00,341.76 779.40,341.76 785.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,330.00 C 771.00,341.76 779.40,341.76 785.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,330.00 C 771.00,341.76 779.40,341.76 785.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,330.00 C 831.00,341.76 839.40,341.76 845.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,330.00 C 831.00,341.76 839.40,341.76 845.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,330.00 C 831.00,341.76 839.40,341.76 845.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,330.00 C 891.00,341.76 899.40,341.76 905.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,330.00 C 891.00,341.76 899.40,341.76 905.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,330.00 C 891.00,341.76 899.40,341.76 905.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,330.00 C 951.00,341.76 959.40,341.76 965.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,330.00 C 951.00,341.76 959.40,341.76 965.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,330.00 C 951.00,341.76 959.40,341.76 965.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,330.00 C 1011.00,341.76 1019.40,341.76 1025.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,330.00 C 1011.00,341.76 1019.40,341.76 1025.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,330.00 C 1011.00,341.76 1019.40,341.76 1025.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,330.00 C 1071.00,341.76 1079.40,341.76 1085.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,330.00 C 1071.00,341.76 1079.40,341.76 1085.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,330.00 C 1071.00,341.76 1079.40,341.76 1085.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,330.00 C 1131.00,341.76 1139.40,341.76 1145.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,330.00 C 1131.00,341.76 1139.40,341.76 1145.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,330.00 C 1131.00,341.76 1139.40,341.76 1145.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,330.00 C 1191.00,341.76 1199.40,341.76 1205.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,330.00 C 1191.00,341.76 1199.40,341.76 1205.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,330.00 C 1191.00,341.76 1199.40,341.76 1205.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,330.00 C 1251.00,341.76 1259.40,341.76 1265.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,330.00 C 1251.00,341.76 1259.40,341.76 1265.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,330.00 C 1251.00,341.76 1259.40,341.76 1265.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,330.00 C 1311.00,341.76 1319.40,341.76 1325.70,330.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,330.00 C 1311.00,341.76 1319.40,341.76 1325.70,330.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,330.00 C 1311.00,341.76 1319.40,341.76 1325.70,330.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,390.00 C 171.00,401.76 179.40,401.76 185.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,390.00 C 171.00,401.76 179.40,401.76 185.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,390.00 C 171.00,401.76 179.40,401.76 185.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,390.00 C 231.00,401.76 239.40,401.76 245.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,390.00 C 231.00,401.76 239.40,401.76 245.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,390.00 C 231.00,401.76 239.40,401.76 245.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,390.00 C 291.00,401.76 299.40,401.76 305.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,390.00 C 291.00,401.76 299.40,401.76 305.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,390.00 C 291.00,401.76 299.40,401.76 305.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,390.00 C 351.00,401.76 359.40,401.76 365.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,390.00 C 351.00,401.76 359.40,401.76 365.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,390.00 C 351.00,401.76 359.40,401.76 365.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,390.00 C 411.00,401.76 419.40,401.76 425.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,390.00 C 411.00,401.76 419.40,401.76 425.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,390.00 C 411.00,401.76 419.40,401.76 425.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,390.00 C 471.00,401.76 479.40,401.76 485.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,390.00 C 471.00,401.76 479.40,401.76 485.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,390.00 C 471.00,401.76 479.40,401.76 485.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,390.00 C 531.00,401.76 539.40,401.76 545.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,390.00 C 531.00,401.76 539.40,401.76 545.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,390.00 C 531.00,401.76 539.40,401.76 545.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,390.00 C 591.00,401.76 599.40,401.76 605.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,390.00 C 591.00,401.76 599.40,401.76 605.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,390.00 C 591.00,401.76 599.40,401.76 605.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,390.00 C 651.00,401.76 659.40,401.76 665.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,390.00 C 651.00,401.76 659.40,401.76 665.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,390.00 C 651.00,401.76 659.40,401.76 665.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,390.00 C 711.00,401.76 719.40,401.76 725.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,390.00 C 711.00,401.76 719.40,401.76 725.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,390.00 C 711.00,401.76 719.40,401.76 725.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,390.00 C 771.00,401.76 779.40,401.76 785.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,390.00 C 771.00,401.76 779.40,401.76 785.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,390.00 C 771.00,401.76 779.40,401.76 785.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,390.00 C 831.00,401.76 839.40,401.76 845.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,390.00 C 831.00,401.76 839.40,401.76 845.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,390.00 C 831.00,401.76 839.40,401.76 845.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,390.00 C 891.00,401.76 899.40,401.76 905.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,390.00 C 891.00,401.76 899.40,401.76 905.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,390.00 C 891.00,401.76 899.40,401.76 905.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,390.00 C 951.00,401.76 959.40,401.76 965.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,390.00 C 951.00,401.76 959.40,401.76 965.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,390.00 C 951.00,401.76 959.40,401.76 965.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,390.00 C 1011.00,401.76 1019.40,401.76 1025.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,390.00 C 1011.00,401.76 1019.40,401.76 1025.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,390.00 C 1011.00,401.76 1019.40,401.76 1025.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,390.00 C 1071.00,401.76 1079.40,401.76 1085.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,390.00 C 1071.00,401.76 1079.40,401.76 1085.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,390.00 C 1071.00,401.76 1079.40,401.76 1085.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,390.00 C 1131.00,401.76 1139.40,401.76 1145.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,390.00 C 1131.00,401.76 1139.40,401.76 1145.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,390.00 C 1131.00,401.76 1139.40,401.76 1145.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,390.00 C 1191.00,401.76 1199.40,401.76 1205.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,390.00 C 1191.00,401.76 1199.40,401.76 1205.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,390.00 C 1191.00,401.76 1199.40,401.76 1205.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,390.00 C 1251.00,401.76 1259.40,401.76 1265.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,390.00 C 1251.00,401.76 1259.40,401.76 1265.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,390.00 C 1251.00,401.76 1259.40,401.76 1265.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,390.00 C 1311.00,401.76 1319.40,401.76 1325.70,390.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,390.00 C 1311.00,401.76 1319.40,401.76 1325.70,390.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,390.00 C 1311.00,401.76 1319.40,401.76 1325.70,390.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,450.00 C 171.00,461.76 179.40,461.76 185.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,450.00 C 171.00,461.76 179.40,461.76 185.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,450.00 C 171.00,461.76 179.40,461.76 185.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,450.00 C 231.00,461.76 239.40,461.76 245.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,450.00 C 231.00,461.76 239.40,461.76 245.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,450.00 C 231.00,461.76 239.40,461.76 245.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,450.00 C 291.00,461.76 299.40,461.76 305.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,450.00 C 291.00,461.76 299.40,461.76 305.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,450.00 C 291.00,461.76 299.40,461.76 305.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,450.00 C 351.00,461.76 359.40,461.76 365.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,450.00 C 351.00,461.76 359.40,461.76 365.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,450.00 C 351.00,461.76 359.40,461.76 365.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,450.00 C 411.00,461.76 419.40,461.76 425.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,450.00 C 411.00,461.76 419.40,461.76 425.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,450.00 C 411.00,461.76 419.40,461.76 425.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,450.00 C 471.00,461.76 479.40,461.76 485.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,450.00 C 471.00,461.76 479.40,461.76 485.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,450.00 C 471.00,461.76 479.40,461.76 485.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,450.00 C 531.00,461.76 539.40,461.76 545.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,450.00 C 531.00,461.76 539.40,461.76 545.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,450.00 C 531.00,461.76 539.40,461.76 545.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,450.00 C 591.00,461.76 599.40,461.76 605.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,450.00 C 591.00,461.76 599.40,461.76 605.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,450.00 C 591.00,461.76 599.40,461.76 605.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,450.00 C 651.00,461.76 659.40,461.76 665.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,450.00 C 651.00,461.76 659.40,461.76 665.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,450.00 C 651.00,461.76 659.40,461.76 665.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,450.00 C 711.00,461.76 719.40,461.76 725.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,450.00 C 711.00,461.76 719.40,461.76 725.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,450.00 C 711.00,461.76 719.40,461.76 725.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,450.00 C 771.00,461.76 779.40,461.76 785.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,450.00 C 771.00,461.76 779.40,461.76 785.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,450.00 C 771.00,461.76 779.40,461.76 785.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,450.00 C 831.00,461.76 839.40,461.76 845.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,450.00 C 831.00,461.76 839.40,461.76 845.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,450.00 C 831.00,461.76 839.40,461.76 845.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,450.00 C 891.00,461.76 899.40,461.76 905.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,450.00 C 891.00,461.76 899.40,461.76 905.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,450.00 C 891.00,461.76 899.40,461.76 905.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,450.00 C 951.00,461.76 959.40,461.76 965.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,450.00 C 951.00,461.76 959.40,461.76 965.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,450.00 C 951.00,461.76 959.40,461.76 965.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,450.00 C 1011.00,461.76 1019.40,461.76 1025.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,450.00 C 1011.00,461.76 1019.40,461.76 1025.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,450.00 C 1011.00,461.76 1019.40,461.76 1025.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,450.00 C 1071.00,461.76 1079.40,461.76 1085.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,450.00 C 1071.00,461.76 1079.40,461.76 1085.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,450.00 C 1071.00,461.76 1079.40,461.76 1085.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,450.00 C 1131.00,461.76 1139.40,461.76 1145.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,450.00 C 1131.00,461.76 1139.40,461.76 1145.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,450.00 C 1131.00,461.76 1139.40,461.76 1145.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,450.00 C 1191.00,461.76 1199.40,461.76 1205.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,450.00 C 1191.00,461.76 1199.40,461.76 1205.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,450.00 C 1191.00,461.76 1199.40,461.76 1205.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,450.00 C 1251.00,461.76 1259.40,461.76 1265.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,450.00 C 1251.00,461.76 1259.40,461.76 1265.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,450.00 C 1251.00,461.76 1259.40,461.76 1265.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,450.00 C 1311.00,461.76 1319.40,461.76 1325.70,450.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,450.00 C 1311.00,461.76 1319.40,461.76 1325.70,450.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,450.00 C 1311.00,461.76 1319.40,461.76 1325.70,450.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,510.00 C 171.00,521.76 179.40,521.76 185.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,510.00 C 171.00,521.76 179.40,521.76 185.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,510.00 C 171.00,521.76 179.40,521.76 185.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,510.00 C 231.00,521.76 239.40,521.76 245.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,510.00 C 231.00,521.76 239.40,521.76 245.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,510.00 C 231.00,521.76 239.40,521.76 245.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,510.00 C 291.00,521.76 299.40,521.76 305.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,510.00 C 291.00,521.76 299.40,521.76 305.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,510.00 C 291.00,521.76 299.40,521.76 305.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,510.00 C 351.00,521.76 359.40,521.76 365.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,510.00 C 351.00,521.76 359.40,521.76 365.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,510.00 C 351.00,521.76 359.40,521.76 365.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,510.00 C 411.00,521.76 419.40,521.76 425.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,510.00 C 411.00,521.76 419.40,521.76 425.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,510.00 C 411.00,521.76 419.40,521.76 425.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,510.00 C 471.00,521.76 479.40,521.76 485.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,510.00 C 471.00,521.76 479.40,521.76 485.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,510.00 C 471.00,521.76 479.40,521.76 485.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,510.00 C 531.00,521.76 539.40,521.76 545.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,510.00 C 531.00,521.76 539.40,521.76 545.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,510.00 C 531.00,521.76 539.40,521.76 545.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,510.00 C 591.00,521.76 599.40,521.76 605.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,510.00 C 591.00,521.76 599.40,521.76 605.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,510.00 C 591.00,521.76 599.40,521.76 605.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,510.00 C 651.00,521.76 659.40,521.76 665.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,510.00 C 651.00,521.76 659.40,521.76 665.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,510.00 C 651.00,521.76 659.40,521.76 665.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,510.00 C 711.00,521.76 719.40,521.76 725.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,510.00 C 711.00,521.76 719.40,521.76 725.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,510.00 C 711.00,521.76 719.40,521.76 725.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,510.00 C 771.00,521.76 779.40,521.76 785.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,510.00 C 771.00,521.76 779.40,521.76 785.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,510.00 C 771.00,521.76 779.40,521.76 785.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,510.00 C 831.00,521.76 839.40,521.76 845.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,510.00 C 831.00,521.76 839.40,521.76 845.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,510.00 C 831.00,521.76 839.40,521.76 845.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,510.00 C 891.00,521.76 899.40,521.76 905.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,510.00 C 891.00,521.76 899.40,521.76 905.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,510.00 C 891.00,521.76 899.40,521.76 905.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,510.00 C 951.00,521.76 959.40,521.76 965.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,510.00 C 951.00,521.76 959.40,521.76 965.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,510.00 C 951.00,521.76 959.40,521.76 965.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,510.00 C 1011.00,521.76 1019.40,521.76 1025.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,510.00 C 1011.00,521.76 1019.40,521.76 1025.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,510.00 C 1011.00,521.76 1019.40,521.76 1025.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,510.00 C 1071.00,521.76 1079.40,521.76 1085.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,510.00 C 1071.00,521.76 1079.40,521.76 1085.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,510.00 C 1071.00,521.76 1079.40,521.76 1085.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,510.00 C 1131.00,521.76 1139.40,521.76 1145.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,510.00 C 1131.00,521.76 1139.40,521.76 1145.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,510.00 C 1131.00,521.76 1139.40,521.76 1145.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,510.00 C 1191.00,521.76 1199.40,521.76 1205.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,510.00 C 1191.00,521.76 1199.40,521.76 1205.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,510.00 C 1191.00,521.76 1199.40,521.76 1205.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,510.00 C 1251.00,521.76 1259.40,521.76 1265.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,510.00 C 1251.00,521.76 1259.40,521.76 1265.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,510.00 C 1251.00,521.76 1259.40,521.76 1265.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,510.00 C 1311.00,521.76 1319.40,521.76 1325.70,510.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,510.00 C 1311.00,521.76 1319.40,521.76 1325.70,510.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,510.00 C 1311.00,521.76 1319.40,521.76 1325.70,510.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,570.00 C 171.00,581.76 179.40,581.76 185.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,570.00 C 171.00,581.76 179.40,581.76 185.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,570.00 C 171.00,581.76 179.40,581.76 185.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,570.00 C 231.00,581.76 239.40,581.76 245.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,570.00 C 231.00,581.76 239.40,581.76 245.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,570.00 C 231.00,581.76 239.40,581.76 245.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,570.00 C 291.00,581.76 299.40,581.76 305.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,570.00 C 291.00,581.76 299.40,581.76 305.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,570.00 C 291.00,581.76 299.40,581.76 305.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,570.00 C 351.00,581.76 359.40,581.76 365.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,570.00 C 351.00,581.76 359.40,581.76 365.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,570.00 C 351.00,581.76 359.40,581.76 365.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,570.00 C 411.00,581.76 419.40,581.76 425.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,570.00 C 411.00,581.76 419.40,581.76 425.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,570.00 C 411.00,581.76 419.40,581.76 425.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,570.00 C 471.00,581.76 479.40,581.76 485.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,570.00 C 471.00,581.76 479.40,581.76 485.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,570.00 C 471.00,581.76 479.40,581.76 485.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,570.00 C 531.00,581.76 539.40,581.76 545.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,570.00 C 531.00,581.76 539.40,581.76 545.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,570.00 C 531.00,581.76 539.40,581.76 545.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,570.00 C 591.00,581.76 599.40,581.76 605.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,570.00 C 591.00,581.76 599.40,581.76 605.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,570.00 C 591.00,581.76 599.40,581.76 605.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,570.00 C 651.00,581.76 659.40,581.76 665.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,570.00 C 651.00,581.76 659.40,581.76 665.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,570.00 C 651.00,581.76 659.40,581.76 665.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,570.00 C 711.00,581.76 719.40,581.76 725.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,570.00 C 711.00,581.76 719.40,581.76 725.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,570.00 C 711.00,581.76 719.40,581.76 725.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,570.00 C 771.00,581.76 779.40,581.76 785.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,570.00 C 771.00,581.76 779.40,581.76 785.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,570.00 C 771.00,581.76 779.40,581.76 785.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,570.00 C 831.00,581.76 839.40,581.76 845.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,570.00 C 831.00,581.76 839.40,581.76 845.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,570.00 C 831.00,581.76 839.40,581.76 845.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,570.00 C 891.00,581.76 899.40,581.76 905.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,570.00 C 891.00,581.76 899.40,581.76 905.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,570.00 C 891.00,581.76 899.40,581.76 905.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,570.00 C 951.00,581.76 959.40,581.76 965.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,570.00 C 951.00,581.76 959.40,581.76 965.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,570.00 C 951.00,581.76 959.40,581.76 965.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,570.00 C 1011.00,581.76 1019.40,581.76 1025.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,570.00 C 1011.00,581.76 1019.40,581.76 1025.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,570.00 C 1011.00,581.76 1019.40,581.76 1025.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,570.00 C 1071.00,581.76 1079.40,581.76 1085.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,570.00 C 1071.00,581.76 1079.40,581.76 1085.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,570.00 C 1071.00,581.76 1079.40,581.76 1085.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,570.00 C 1131.00,581.76 1139.40,581.76 1145.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,570.00 C 1131.00,581.76 1139.40,581.76 1145.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,570.00 C 1131.00,581.76 1139.40,581.76 1145.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,570.00 C 1191.00,581.76 1199.40,581.76 1205.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,570.00 C 1191.00,581.76 1199.40,581.76 1205.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,570.00 C 1191.00,581.76 1199.40,581.76 1205.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,570.00 C 1251.00,581.76 1259.40,581.76 1265.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,570.00 C 1251.00,581.76 1259.40,581.76 1265.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,570.00 C 1251.00,581.76 1259.40,581.76 1265.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,570.00 C 1311.00,581.76 1319.40,581.76 1325.70,570.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,570.00 C 1311.00,581.76 1319.40,581.76 1325.70,570.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,570.00 C 1311.00,581.76 1319.40,581.76 1325.70,570.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,630.00 C 171.00,641.76 179.40,641.76 185.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,630.00 C 171.00,641.76 179.40,641.76 185.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,630.00 C 171.00,641.76 179.40,641.76 185.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,630.00 C 231.00,641.76 239.40,641.76 245.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,630.00 C 231.00,641.76 239.40,641.76 245.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,630.00 C 231.00,641.76 239.40,641.76 245.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,630.00 C 291.00,641.76 299.40,641.76 305.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,630.00 C 291.00,641.76 299.40,641.76 305.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,630.00 C 291.00,641.76 299.40,641.76 305.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,630.00 C 351.00,641.76 359.40,641.76 365.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,630.00 C 351.00,641.76 359.40,641.76 365.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,630.00 C 351.00,641.76 359.40,641.76 365.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,630.00 C 411.00,641.76 419.40,641.76 425.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,630.00 C 411.00,641.76 419.40,641.76 425.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,630.00 C 411.00,641.76 419.40,641.76 425.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,630.00 C 471.00,641.76 479.40,641.76 485.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,630.00 C 471.00,641.76 479.40,641.76 485.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,630.00 C 471.00,641.76 479.40,641.76 485.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,630.00 C 531.00,641.76 539.40,641.76 545.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,630.00 C 531.00,641.76 539.40,641.76 545.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,630.00 C 531.00,641.76 539.40,641.76 545.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,630.00 C 591.00,641.76 599.40,641.76 605.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,630.00 C 591.00,641.76 599.40,641.76 605.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,630.00 C 591.00,641.76 599.40,641.76 605.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,630.00 C 651.00,641.76 659.40,641.76 665.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,630.00 C 651.00,641.76 659.40,641.76 665.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,630.00 C 651.00,641.76 659.40,641.76 665.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,630.00 C 711.00,641.76 719.40,641.76 725.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,630.00 C 711.00,641.76 719.40,641.76 725.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,630.00 C 711.00,641.76 719.40,641.76 725.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,630.00 C 771.00,641.76 779.40,641.76 785.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,630.00 C 771.00,641.76 779.40,641.76 785.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,630.00 C 771.00,641.76 779.40,641.76 785.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,630.00 C 831.00,641.76 839.40,641.76 845.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,630.00 C 831.00,641.76 839.40,641.76 845.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,630.00 C 831.00,641.76 839.40,641.76 845.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,630.00 C 891.00,641.76 899.40,641.76 905.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,630.00 C 891.00,641.76 899.40,641.76 905.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,630.00 C 891.00,641.76 899.40,641.76 905.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,630.00 C 951.00,641.76 959.40,641.76 965.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,630.00 C 951.00,641.76 959.40,641.76 965.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,630.00 C 951.00,641.76 959.40,641.76 965.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,630.00 C 1011.00,641.76 1019.40,641.76 1025.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,630.00 C 1011.00,641.76 1019.40,641.76 1025.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,630.00 C 1011.00,641.76 1019.40,641.76 1025.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,630.00 C 1071.00,641.76 1079.40,641.76 1085.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,630.00 C 1071.00,641.76 1079.40,641.76 1085.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,630.00 C 1071.00,641.76 1079.40,641.76 1085.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,630.00 C 1131.00,641.76 1139.40,641.76 1145.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,630.00 C 1131.00,641.76 1139.40,641.76 1145.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,630.00 C 1131.00,641.76 1139.40,641.76 1145.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,630.00 C 1191.00,641.76 1199.40,641.76 1205.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,630.00 C 1191.00,641.76 1199.40,641.76 1205.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,630.00 C 1191.00,641.76 1199.40,641.76 1205.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,630.00 C 1251.00,641.76 1259.40,641.76 1265.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,630.00 C 1251.00,641.76 1259.40,641.76 1265.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,630.00 C 1251.00,641.76 1259.40,641.76 1265.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,630.00 C 1311.00,641.76 1319.40,641.76 1325.70,630.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,630.00 C 1311.00,641.76 1319.40,641.76 1325.70,630.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,630.00 C 1311.00,641.76 1319.40,641.76 1325.70,630.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,690.00 C 171.00,701.76 179.40,701.76 185.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,690.00 C 171.00,701.76 179.40,701.76 185.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,690.00 C 171.00,701.76 179.40,701.76 185.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,690.00 C 231.00,701.76 239.40,701.76 245.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,690.00 C 231.00,701.76 239.40,701.76 245.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,690.00 C 231.00,701.76 239.40,701.76 245.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,690.00 C 291.00,701.76 299.40,701.76 305.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,690.00 C 291.00,701.76 299.40,701.76 305.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,690.00 C 291.00,701.76 299.40,701.76 305.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,690.00 C 351.00,701.76 359.40,701.76 365.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,690.00 C 351.00,701.76 359.40,701.76 365.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,690.00 C 351.00,701.76 359.40,701.76 365.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,690.00 C 411.00,701.76 419.40,701.76 425.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,690.00 C 411.00,701.76 419.40,701.76 425.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,690.00 C 411.00,701.76 419.40,701.76 425.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,690.00 C 471.00,701.76 479.40,701.76 485.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,690.00 C 471.00,701.76 479.40,701.76 485.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,690.00 C 471.00,701.76 479.40,701.76 485.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,690.00 C 531.00,701.76 539.40,701.76 545.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,690.00 C 531.00,701.76 539.40,701.76 545.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,690.00 C 531.00,701.76 539.40,701.76 545.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,690.00 C 591.00,701.76 599.40,701.76 605.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,690.00 C 591.00,701.76 599.40,701.76 605.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,690.00 C 591.00,701.76 599.40,701.76 605.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,690.00 C 651.00,701.76 659.40,701.76 665.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,690.00 C 651.00,701.76 659.40,701.76 665.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,690.00 C 651.00,701.76 659.40,701.76 665.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,690.00 C 711.00,701.76 719.40,701.76 725.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,690.00 C 711.00,701.76 719.40,701.76 725.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,690.00 C 711.00,701.76 719.40,701.76 725.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,690.00 C 771.00,701.76 779.40,701.76 785.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,690.00 C 771.00,701.76 779.40,701.76 785.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,690.00 C 771.00,701.76 779.40,701.76 785.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,690.00 C 831.00,701.76 839.40,701.76 845.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,690.00 C 831.00,701.76 839.40,701.76 845.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,690.00 C 831.00,701.76 839.40,701.76 845.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,690.00 C 891.00,701.76 899.40,701.76 905.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,690.00 C 891.00,701.76 899.40,701.76 905.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,690.00 C 891.00,701.76 899.40,701.76 905.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,690.00 C 951.00,701.76 959.40,701.76 965.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,690.00 C 951.00,701.76 959.40,701.76 965.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,690.00 C 951.00,701.76 959.40,701.76 965.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,690.00 C 1011.00,701.76 1019.40,701.76 1025.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,690.00 C 1011.00,701.76 1019.40,701.76 1025.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,690.00 C 1011.00,701.76 1019.40,701.76 1025.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,690.00 C 1071.00,701.76 1079.40,701.76 1085.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,690.00 C 1071.00,701.76 1079.40,701.76 1085.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,690.00 C 1071.00,701.76 1079.40,701.76 1085.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,690.00 C 1131.00,701.76 1139.40,701.76 1145.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,690.00 C 1131.00,701.76 1139.40,701.76 1145.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,690.00 C 1131.00,701.76 1139.40,701.76 1145.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,690.00 C 1191.00,701.76 1199.40,701.76 1205.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,690.00 C 1191.00,701.76 1199.40,701.76 1205.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,690.00 C 1191.00,701.76 1199.40,701.76 1205.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,690.00 C 1251.00,701.76 1259.40,701.76 1265.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,690.00 C 1251.00,701.76 1259.40,701.76 1265.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,690.00 C 1251.00,701.76 1259.40,701.76 1265.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,690.00 C 1311.00,701.76 1319.40,701.76 1325.70,690.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,690.00 C 1311.00,701.76 1319.40,701.76 1325.70,690.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,690.00 C 1311.00,701.76 1319.40,701.76 1325.70,690.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,750.00 C 171.00,761.76 179.40,761.76 185.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,750.00 C 171.00,761.76 179.40,761.76 185.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,750.00 C 171.00,761.76 179.40,761.76 185.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,750.00 C 231.00,761.76 239.40,761.76 245.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,750.00 C 231.00,761.76 239.40,761.76 245.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,750.00 C 231.00,761.76 239.40,761.76 245.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,750.00 C 291.00,761.76 299.40,761.76 305.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,750.00 C 291.00,761.76 299.40,761.76 305.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,750.00 C 291.00,761.76 299.40,761.76 305.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,750.00 C 351.00,761.76 359.40,761.76 365.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,750.00 C 351.00,761.76 359.40,761.76 365.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,750.00 C 351.00,761.76 359.40,761.76 365.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,750.00 C 411.00,761.76 419.40,761.76 425.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,750.00 C 411.00,761.76 419.40,761.76 425.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,750.00 C 411.00,761.76 419.40,761.76 425.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,750.00 C 471.00,761.76 479.40,761.76 485.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,750.00 C 471.00,761.76 479.40,761.76 485.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,750.00 C 471.00,761.76 479.40,761.76 485.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,750.00 C 531.00,761.76 539.40,761.76 545.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,750.00 C 531.00,761.76 539.40,761.76 545.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,750.00 C 531.00,761.76 539.40,761.76 545.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,750.00 C 591.00,761.76 599.40,761.76 605.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,750.00 C 591.00,761.76 599.40,761.76 605.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,750.00 C 591.00,761.76 599.40,761.76 605.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,750.00 C 651.00,761.76 659.40,761.76 665.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,750.00 C 651.00,761.76 659.40,761.76 665.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,750.00 C 651.00,761.76 659.40,761.76 665.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,750.00 C 711.00,761.76 719.40,761.76 725.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,750.00 C 711.00,761.76 719.40,761.76 725.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,750.00 C 711.00,761.76 719.40,761.76 725.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,750.00 C 771.00,761.76 779.40,761.76 785.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,750.00 C 771.00,761.76 779.40,761.76 785.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,750.00 C 771.00,761.76 779.40,761.76 785.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,750.00 C 831.00,761.76 839.40,761.76 845.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,750.00 C 831.00,761.76 839.40,761.76 845.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,750.00 C 831.00,761.76 839.40,761.76 845.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,750.00 C 891.00,761.76 899.40,761.76 905.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,750.00 C 891.00,761.76 899.40,761.76 905.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,750.00 C 891.00,761.76 899.40,761.76 905.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,750.00 C 951.00,761.76 959.40,761.76 965.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,750.00 C 951.00,761.76 959.40,761.76 965.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,750.00 C 951.00,761.76 959.40,761.76 965.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,750.00 C 1011.00,761.76 1019.40,761.76 1025.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,750.00 C 1011.00,761.76 1019.40,761.76 1025.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,750.00 C 1011.00,761.76 1019.40,761.76 1025.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,750.00 C 1071.00,761.76 1079.40,761.76 1085.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,750.00 C 1071.00,761.76 1079.40,761.76 1085.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,750.00 C 1071.00,761.76 1079.40,761.76 1085.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,750.00 C 1131.00,761.76 1139.40,761.76 1145.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,750.00 C 1131.00,761.76 1139.40,761.76 1145.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,750.00 C 1131.00,761.76 1139.40,761.76 1145.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,750.00 C 1191.00,761.76 1199.40,761.76 1205.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,750.00 C 1191.00,761.76 1199.40,761.76 1205.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,750.00 C 1191.00,761.76 1199.40,761.76 1205.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,750.00 C 1251.00,761.76 1259.40,761.76 1265.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,750.00 C 1251.00,761.76 1259.40,761.76 1265.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,750.00 C 1251.00,761.76 1259.40,761.76 1265.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,750.00 C 1311.00,761.76 1319.40,761.76 1325.70,750.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,750.00 C 1311.00,761.76 1319.40,761.76 1325.70,750.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,750.00 C 1311.00,761.76 1319.40,761.76 1325.70,750.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,810.00 C 171.00,821.76 179.40,821.76 185.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,810.00 C 171.00,821.76 179.40,821.76 185.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,810.00 C 171.00,821.76 179.40,821.76 185.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,810.00 C 231.00,821.76 239.40,821.76 245.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,810.00 C 231.00,821.76 239.40,821.76 245.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,810.00 C 231.00,821.76 239.40,821.76 245.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,810.00 C 291.00,821.76 299.40,821.76 305.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,810.00 C 291.00,821.76 299.40,821.76 305.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,810.00 C 291.00,821.76 299.40,821.76 305.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,810.00 C 351.00,821.76 359.40,821.76 365.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,810.00 C 351.00,821.76 359.40,821.76 365.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,810.00 C 351.00,821.76 359.40,821.76 365.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,810.00 C 411.00,821.76 419.40,821.76 425.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,810.00 C 411.00,821.76 419.40,821.76 425.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,810.00 C 411.00,821.76 419.40,821.76 425.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,810.00 C 471.00,821.76 479.40,821.76 485.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,810.00 C 471.00,821.76 479.40,821.76 485.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,810.00 C 471.00,821.76 479.40,821.76 485.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,810.00 C 531.00,821.76 539.40,821.76 545.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,810.00 C 531.00,821.76 539.40,821.76 545.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,810.00 C 531.00,821.76 539.40,821.76 545.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,810.00 C 591.00,821.76 599.40,821.76 605.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,810.00 C 591.00,821.76 599.40,821.76 605.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,810.00 C 591.00,821.76 599.40,821.76 605.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,810.00 C 651.00,821.76 659.40,821.76 665.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,810.00 C 651.00,821.76 659.40,821.76 665.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,810.00 C 651.00,821.76 659.40,821.76 665.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,810.00 C 711.00,821.76 719.40,821.76 725.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,810.00 C 711.00,821.76 719.40,821.76 725.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,810.00 C 711.00,821.76 719.40,821.76 725.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,810.00 C 771.00,821.76 779.40,821.76 785.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,810.00 C 771.00,821.76 779.40,821.76 785.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,810.00 C 771.00,821.76 779.40,821.76 785.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,810.00 C 831.00,821.76 839.40,821.76 845.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,810.00 C 831.00,821.76 839.40,821.76 845.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,810.00 C 831.00,821.76 839.40,821.76 845.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,810.00 C 891.00,821.76 899.40,821.76 905.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,810.00 C 891.00,821.76 899.40,821.76 905.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,810.00 C 891.00,821.76 899.40,821.76 905.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,810.00 C 951.00,821.76 959.40,821.76 965.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,810.00 C 951.00,821.76 959.40,821.76 965.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,810.00 C 951.00,821.76 959.40,821.76 965.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,810.00 C 1011.00,821.76 1019.40,821.76 1025.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,810.00 C 1011.00,821.76 1019.40,821.76 1025.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,810.00 C 1011.00,821.76 1019.40,821.76 1025.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,810.00 C 1071.00,821.76 1079.40,821.76 1085.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,810.00 C 1071.00,821.76 1079.40,821.76 1085.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,810.00 C 1071.00,821.76 1079.40,821.76 1085.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,810.00 C 1131.00,821.76 1139.40,821.76 1145.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,810.00 C 1131.00,821.76 1139.40,821.76 1145.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,810.00 C 1131.00,821.76 1139.40,821.76 1145.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,810.00 C 1191.00,821.76 1199.40,821.76 1205.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,810.00 C 1191.00,821.76 1199.40,821.76 1205.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,810.00 C 1191.00,821.76 1199.40,821.76 1205.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,810.00 C 1251.00,821.76 1259.40,821.76 1265.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,810.00 C 1251.00,821.76 1259.40,821.76 1265.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,810.00 C 1251.00,821.76 1259.40,821.76 1265.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,810.00 C 1311.00,821.76 1319.40,821.76 1325.70,810.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,810.00 C 1311.00,821.76 1319.40,821.76 1325.70,810.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,810.00 C 1311.00,821.76 1319.40,821.76 1325.70,810.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,870.00 C 171.00,881.76 179.40,881.76 185.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,870.00 C 171.00,881.76 179.40,881.76 185.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,870.00 C 171.00,881.76 179.40,881.76 185.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,870.00 C 231.00,881.76 239.40,881.76 245.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,870.00 C 231.00,881.76 239.40,881.76 245.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,870.00 C 231.00,881.76 239.40,881.76 245.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,870.00 C 291.00,881.76 299.40,881.76 305.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,870.00 C 291.00,881.76 299.40,881.76 305.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,870.00 C 291.00,881.76 299.40,881.76 305.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,870.00 C 351.00,881.76 359.40,881.76 365.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,870.00 C 351.00,881.76 359.40,881.76 365.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,870.00 C 351.00,881.76 359.40,881.76 365.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,870.00 C 411.00,881.76 419.40,881.76 425.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,870.00 C 411.00,881.76 419.40,881.76 425.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,870.00 C 411.00,881.76 419.40,881.76 425.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,870.00 C 471.00,881.76 479.40,881.76 485.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,870.00 C 471.00,881.76 479.40,881.76 485.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,870.00 C 471.00,881.76 479.40,881.76 485.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,870.00 C 531.00,881.76 539.40,881.76 545.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,870.00 C 531.00,881.76 539.40,881.76 545.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,870.00 C 531.00,881.76 539.40,881.76 545.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,870.00 C 591.00,881.76 599.40,881.76 605.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,870.00 C 591.00,881.76 599.40,881.76 605.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,870.00 C 591.00,881.76 599.40,881.76 605.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,870.00 C 651.00,881.76 659.40,881.76 665.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,870.00 C 651.00,881.76 659.40,881.76 665.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,870.00 C 651.00,881.76 659.40,881.76 665.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,870.00 C 711.00,881.76 719.40,881.76 725.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,870.00 C 711.00,881.76 719.40,881.76 725.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,870.00 C 711.00,881.76 719.40,881.76 725.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,870.00 C 771.00,881.76 779.40,881.76 785.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,870.00 C 771.00,881.76 779.40,881.76 785.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,870.00 C 771.00,881.76 779.40,881.76 785.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,870.00 C 831.00,881.76 839.40,881.76 845.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,870.00 C 831.00,881.76 839.40,881.76 845.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,870.00 C 831.00,881.76 839.40,881.76 845.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,870.00 C 891.00,881.76 899.40,881.76 905.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,870.00 C 891.00,881.76 899.40,881.76 905.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,870.00 C 891.00,881.76 899.40,881.76 905.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,870.00 C 951.00,881.76 959.40,881.76 965.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,870.00 C 951.00,881.76 959.40,881.76 965.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,870.00 C 951.00,881.76 959.40,881.76 965.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,870.00 C 1011.00,881.76 1019.40,881.76 1025.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,870.00 C 1011.00,881.76 1019.40,881.76 1025.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,870.00 C 1011.00,881.76 1019.40,881.76 1025.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,870.00 C 1071.00,881.76 1079.40,881.76 1085.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,870.00 C 1071.00,881.76 1079.40,881.76 1085.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,870.00 C 1071.00,881.76 1079.40,881.76 1085.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,870.00 C 1131.00,881.76 1139.40,881.76 1145.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,870.00 C 1131.00,881.76 1139.40,881.76 1145.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,870.00 C 1131.00,881.76 1139.40,881.76 1145.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,870.00 C 1191.00,881.76 1199.40,881.76 1205.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,870.00 C 1191.00,881.76 1199.40,881.76 1205.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,870.00 C 1191.00,881.76 1199.40,881.76 1205.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,870.00 C 1251.00,881.76 1259.40,881.76 1265.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,870.00 C 1251.00,881.76 1259.40,881.76 1265.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,870.00 C 1251.00,881.76 1259.40,881.76 1265.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,870.00 C 1311.00,881.76 1319.40,881.76 1325.70,870.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,870.00 C 1311.00,881.76 1319.40,881.76 1325.70,870.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,870.00 C 1311.00,881.76 1319.40,881.76 1325.70,870.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,930.00 C 171.00,941.76 179.40,941.76 185.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,930.00 C 171.00,941.76 179.40,941.76 185.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,930.00 C 171.00,941.76 179.40,941.76 185.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,930.00 C 231.00,941.76 239.40,941.76 245.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,930.00 C 231.00,941.76 239.40,941.76 245.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,930.00 C 231.00,941.76 239.40,941.76 245.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,930.00 C 291.00,941.76 299.40,941.76 305.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,930.00 C 291.00,941.76 299.40,941.76 305.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,930.00 C 291.00,941.76 299.40,941.76 305.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,930.00 C 351.00,941.76 359.40,941.76 365.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,930.00 C 351.00,941.76 359.40,941.76 365.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,930.00 C 351.00,941.76 359.40,941.76 365.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,930.00 C 411.00,941.76 419.40,941.76 425.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,930.00 C 411.00,941.76 419.40,941.76 425.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,930.00 C 411.00,941.76 419.40,941.76 425.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,930.00 C 471.00,941.76 479.40,941.76 485.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,930.00 C 471.00,941.76 479.40,941.76 485.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,930.00 C 471.00,941.76 479.40,941.76 485.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,930.00 C 531.00,941.76 539.40,941.76 545.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,930.00 C 531.00,941.76 539.40,941.76 545.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,930.00 C 531.00,941.76 539.40,941.76 545.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,930.00 C 591.00,941.76 599.40,941.76 605.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,930.00 C 591.00,941.76 599.40,941.76 605.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,930.00 C 591.00,941.76 599.40,941.76 605.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,930.00 C 651.00,941.76 659.40,941.76 665.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,930.00 C 651.00,941.76 659.40,941.76 665.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,930.00 C 651.00,941.76 659.40,941.76 665.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,930.00 C 711.00,941.76 719.40,941.76 725.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,930.00 C 711.00,941.76 719.40,941.76 725.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,930.00 C 711.00,941.76 719.40,941.76 725.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,930.00 C 771.00,941.76 779.40,941.76 785.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,930.00 C 771.00,941.76 779.40,941.76 785.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,930.00 C 771.00,941.76 779.40,941.76 785.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,930.00 C 831.00,941.76 839.40,941.76 845.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,930.00 C 831.00,941.76 839.40,941.76 845.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,930.00 C 831.00,941.76 839.40,941.76 845.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,930.00 C 891.00,941.76 899.40,941.76 905.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,930.00 C 891.00,941.76 899.40,941.76 905.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,930.00 C 891.00,941.76 899.40,941.76 905.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,930.00 C 951.00,941.76 959.40,941.76 965.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,930.00 C 951.00,941.76 959.40,941.76 965.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,930.00 C 951.00,941.76 959.40,941.76 965.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,930.00 C 1011.00,941.76 1019.40,941.76 1025.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,930.00 C 1011.00,941.76 1019.40,941.76 1025.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,930.00 C 1011.00,941.76 1019.40,941.76 1025.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,930.00 C 1071.00,941.76 1079.40,941.76 1085.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,930.00 C 1071.00,941.76 1079.40,941.76 1085.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,930.00 C 1071.00,941.76 1079.40,941.76 1085.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,930.00 C 1131.00,941.76 1139.40,941.76 1145.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,930.00 C 1131.00,941.76 1139.40,941.76 1145.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,930.00 C 1131.00,941.76 1139.40,941.76 1145.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,930.00 C 1191.00,941.76 1199.40,941.76 1205.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,930.00 C 1191.00,941.76 1199.40,941.76 1205.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,930.00 C 1191.00,941.76 1199.40,941.76 1205.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,930.00 C 1251.00,941.76 1259.40,941.76 1265.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,930.00 C 1251.00,941.76 1259.40,941.76 1265.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,930.00 C 1251.00,941.76 1259.40,941.76 1265.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,930.00 C 1311.00,941.76 1319.40,941.76 1325.70,930.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,930.00 C 1311.00,941.76 1319.40,941.76 1325.70,930.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,930.00 C 1311.00,941.76 1319.40,941.76 1325.70,930.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,990.00 C 171.00,1001.76 179.40,1001.76 185.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,990.00 C 171.00,1001.76 179.40,1001.76 185.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,990.00 C 171.00,1001.76 179.40,1001.76 185.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,990.00 C 231.00,1001.76 239.40,1001.76 245.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,990.00 C 231.00,1001.76 239.40,1001.76 245.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,990.00 C 231.00,1001.76 239.40,1001.76 245.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,990.00 C 291.00,1001.76 299.40,1001.76 305.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,990.00 C 291.00,1001.76 299.40,1001.76 305.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,990.00 C 291.00,1001.76 299.40,1001.76 305.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,990.00 C 351.00,1001.76 359.40,1001.76 365.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,990.00 C 351.00,1001.76 359.40,1001.76 365.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,990.00 C 351.00,1001.76 359.40,1001.76 365.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,990.00 C 411.00,1001.76 419.40,1001.76 425.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,990.00 C 411.00,1001.76 419.40,1001.76 425.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,990.00 C 411.00,1001.76 419.40,1001.76 425.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,990.00 C 471.00,1001.76 479.40,1001.76 485.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,990.00 C 471.00,1001.76 479.40,1001.76 485.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,990.00 C 471.00,1001.76 479.40,1001.76 485.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,990.00 C 531.00,1001.76 539.40,1001.76 545.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,990.00 C 531.00,1001.76 539.40,1001.76 545.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,990.00 C 531.00,1001.76 539.40,1001.76 545.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,990.00 C 591.00,1001.76 599.40,1001.76 605.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,990.00 C 591.00,1001.76 599.40,1001.76 605.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,990.00 C 591.00,1001.76 599.40,1001.76 605.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,990.00 C 651.00,1001.76 659.40,1001.76 665.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,990.00 C 651.00,1001.76 659.40,1001.76 665.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,990.00 C 651.00,1001.76 659.40,1001.76 665.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,990.00 C 711.00,1001.76 719.40,1001.76 725.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,990.00 C 711.00,1001.76 719.40,1001.76 725.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,990.00 C 711.00,1001.76 719.40,1001.76 725.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,990.00 C 771.00,1001.76 779.40,1001.76 785.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,990.00 C 771.00,1001.76 779.40,1001.76 785.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,990.00 C 771.00,1001.76 779.40,1001.76 785.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,990.00 C 831.00,1001.76 839.40,1001.76 845.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,990.00 C 831.00,1001.76 839.40,1001.76 845.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,990.00 C 831.00,1001.76 839.40,1001.76 845.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,990.00 C 891.00,1001.76 899.40,1001.76 905.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,990.00 C 891.00,1001.76 899.40,1001.76 905.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,990.00 C 891.00,1001.76 899.40,1001.76 905.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,990.00 C 951.00,1001.76 959.40,1001.76 965.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,990.00 C 951.00,1001.76 959.40,1001.76 965.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,990.00 C 951.00,1001.76 959.40,1001.76 965.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,990.00 C 1011.00,1001.76 1019.40,1001.76 1025.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,990.00 C 1011.00,1001.76 1019.40,1001.76 1025.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,990.00 C 1011.00,1001.76 1019.40,1001.76 1025.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,990.00 C 1071.00,1001.76 1079.40,1001.76 1085.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,990.00 C 1071.00,1001.76 1079.40,1001.76 1085.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,990.00 C 1071.00,1001.76 1079.40,1001.76 1085.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,990.00 C 1131.00,1001.76 1139.40,1001.76 1145.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,990.00 C 1131.00,1001.76 1139.40,1001.76 1145.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,990.00 C 1131.00,1001.76 1139.40,1001.76 1145.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,990.00 C 1191.00,1001.76 1199.40,1001.76 1205.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,990.00 C 1191.00,1001.76 1199.40,1001.76 1205.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,990.00 C 1191.00,1001.76 1199.40,1001.76 1205.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,990.00 C 1251.00,1001.76 1259.40,1001.76 1265.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,990.00 C 1251.00,1001.76 1259.40,1001.76 1265.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,990.00 C 1251.00,1001.76 1259.40,1001.76 1265.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,990.00 C 1311.00,1001.76 1319.40,1001.76 1325.70,990.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,990.00 C 1311.00,1001.76 1319.40,1001.76 1325.70,990.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,990.00 C 1311.00,1001.76 1319.40,1001.76 1325.70,990.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,1050.00 C 171.00,1061.76 179.40,1061.76 185.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,1050.00 C 171.00,1061.76 179.40,1061.76 185.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,1050.00 C 171.00,1061.76 179.40,1061.76 185.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,1050.00 C 231.00,1061.76 239.40,1061.76 245.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,1050.00 C 231.00,1061.76 239.40,1061.76 245.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,1050.00 C 231.00,1061.76 239.40,1061.76 245.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,1050.00 C 291.00,1061.76 299.40,1061.76 305.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,1050.00 C 291.00,1061.76 299.40,1061.76 305.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,1050.00 C 291.00,1061.76 299.40,1061.76 305.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,1050.00 C 351.00,1061.76 359.40,1061.76 365.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,1050.00 C 351.00,1061.76 359.40,1061.76 365.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,1050.00 C 351.00,1061.76 359.40,1061.76 365.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,1050.00 C 411.00,1061.76 419.40,1061.76 425.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,1050.00 C 411.00,1061.76 419.40,1061.76 425.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,1050.00 C 411.00,1061.76 419.40,1061.76 425.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,1050.00 C 471.00,1061.76 479.40,1061.76 485.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,1050.00 C 471.00,1061.76 479.40,1061.76 485.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,1050.00 C 471.00,1061.76 479.40,1061.76 485.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,1050.00 C 531.00,1061.76 539.40,1061.76 545.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,1050.00 C 531.00,1061.76 539.40,1061.76 545.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,1050.00 C 531.00,1061.76 539.40,1061.76 545.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,1050.00 C 591.00,1061.76 599.40,1061.76 605.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,1050.00 C 591.00,1061.76 599.40,1061.76 605.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,1050.00 C 591.00,1061.76 599.40,1061.76 605.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,1050.00 C 651.00,1061.76 659.40,1061.76 665.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,1050.00 C 651.00,1061.76 659.40,1061.76 665.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,1050.00 C 651.00,1061.76 659.40,1061.76 665.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,1050.00 C 711.00,1061.76 719.40,1061.76 725.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,1050.00 C 711.00,1061.76 719.40,1061.76 725.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,1050.00 C 711.00,1061.76 719.40,1061.76 725.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,1050.00 C 771.00,1061.76 779.40,1061.76 785.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,1050.00 C 771.00,1061.76 779.40,1061.76 785.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,1050.00 C 771.00,1061.76 779.40,1061.76 785.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,1050.00 C 831.00,1061.76 839.40,1061.76 845.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,1050.00 C 831.00,1061.76 839.40,1061.76 845.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,1050.00 C 831.00,1061.76 839.40,1061.76 845.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,1050.00 C 891.00,1061.76 899.40,1061.76 905.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,1050.00 C 891.00,1061.76 899.40,1061.76 905.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,1050.00 C 891.00,1061.76 899.40,1061.76 905.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,1050.00 C 951.00,1061.76 959.40,1061.76 965.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,1050.00 C 951.00,1061.76 959.40,1061.76 965.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,1050.00 C 951.00,1061.76 959.40,1061.76 965.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,1050.00 C 1011.00,1061.76 1019.40,1061.76 1025.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,1050.00 C 1011.00,1061.76 1019.40,1061.76 1025.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,1050.00 C 1011.00,1061.76 1019.40,1061.76 1025.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,1050.00 C 1071.00,1061.76 1079.40,1061.76 1085.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,1050.00 C 1071.00,1061.76 1079.40,1061.76 1085.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,1050.00 C 1071.00,1061.76 1079.40,1061.76 1085.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,1050.00 C 1131.00,1061.76 1139.40,1061.76 1145.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,1050.00 C 1131.00,1061.76 1139.40,1061.76 1145.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,1050.00 C 1131.00,1061.76 1139.40,1061.76 1145.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,1050.00 C 1191.00,1061.76 1199.40,1061.76 1205.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,1050.00 C 1191.00,1061.76 1199.40,1061.76 1205.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,1050.00 C 1191.00,1061.76 1199.40,1061.76 1205.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,1050.00 C 1251.00,1061.76 1259.40,1061.76 1265.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,1050.00 C 1251.00,1061.76 1259.40,1061.76 1265.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,1050.00 C 1251.00,1061.76 1259.40,1061.76 1265.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,1050.00 C 1311.00,1061.76 1319.40,1061.76 1325.70,1050.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,1050.00 C 1311.00,1061.76 1319.40,1061.76 1325.70,1050.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,1050.00 C 1311.00,1061.76 1319.40,1061.76 1325.70,1050.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,1110.00 C 171.00,1121.76 179.40,1121.76 185.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,1110.00 C 171.00,1121.76 179.40,1121.76 185.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,1110.00 C 171.00,1121.76 179.40,1121.76 185.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,1110.00 C 231.00,1121.76 239.40,1121.76 245.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,1110.00 C 231.00,1121.76 239.40,1121.76 245.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,1110.00 C 231.00,1121.76 239.40,1121.76 245.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,1110.00 C 291.00,1121.76 299.40,1121.76 305.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,1110.00 C 291.00,1121.76 299.40,1121.76 305.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,1110.00 C 291.00,1121.76 299.40,1121.76 305.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,1110.00 C 351.00,1121.76 359.40,1121.76 365.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,1110.00 C 351.00,1121.76 359.40,1121.76 365.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,1110.00 C 351.00,1121.76 359.40,1121.76 365.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,1110.00 C 411.00,1121.76 419.40,1121.76 425.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,1110.00 C 411.00,1121.76 419.40,1121.76 425.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,1110.00 C 411.00,1121.76 419.40,1121.76 425.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,1110.00 C 471.00,1121.76 479.40,1121.76 485.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,1110.00 C 471.00,1121.76 479.40,1121.76 485.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,1110.00 C 471.00,1121.76 479.40,1121.76 485.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,1110.00 C 531.00,1121.76 539.40,1121.76 545.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,1110.00 C 531.00,1121.76 539.40,1121.76 545.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,1110.00 C 531.00,1121.76 539.40,1121.76 545.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,1110.00 C 591.00,1121.76 599.40,1121.76 605.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,1110.00 C 591.00,1121.76 599.40,1121.76 605.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,1110.00 C 591.00,1121.76 599.40,1121.76 605.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,1110.00 C 651.00,1121.76 659.40,1121.76 665.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,1110.00 C 651.00,1121.76 659.40,1121.76 665.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,1110.00 C 651.00,1121.76 659.40,1121.76 665.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,1110.00 C 711.00,1121.76 719.40,1121.76 725.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,1110.00 C 711.00,1121.76 719.40,1121.76 725.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,1110.00 C 711.00,1121.76 719.40,1121.76 725.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,1110.00 C 771.00,1121.76 779.40,1121.76 785.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,1110.00 C 771.00,1121.76 779.40,1121.76 785.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,1110.00 C 771.00,1121.76 779.40,1121.76 785.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,1110.00 C 831.00,1121.76 839.40,1121.76 845.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,1110.00 C 831.00,1121.76 839.40,1121.76 845.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,1110.00 C 831.00,1121.76 839.40,1121.76 845.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,1110.00 C 891.00,1121.76 899.40,1121.76 905.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,1110.00 C 891.00,1121.76 899.40,1121.76 905.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,1110.00 C 891.00,1121.76 899.40,1121.76 905.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,1110.00 C 951.00,1121.76 959.40,1121.76 965.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,1110.00 C 951.00,1121.76 959.40,1121.76 965.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,1110.00 C 951.00,1121.76 959.40,1121.76 965.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,1110.00 C 1011.00,1121.76 1019.40,1121.76 1025.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,1110.00 C 1011.00,1121.76 1019.40,1121.76 1025.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,1110.00 C 1011.00,1121.76 1019.40,1121.76 1025.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,1110.00 C 1071.00,1121.76 1079.40,1121.76 1085.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,1110.00 C 1071.00,1121.76 1079.40,1121.76 1085.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,1110.00 C 1071.00,1121.76 1079.40,1121.76 1085.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,1110.00 C 1131.00,1121.76 1139.40,1121.76 1145.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,1110.00 C 1131.00,1121.76 1139.40,1121.76 1145.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,1110.00 C 1131.00,1121.76 1139.40,1121.76 1145.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,1110.00 C 1191.00,1121.76 1199.40,1121.76 1205.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,1110.00 C 1191.00,1121.76 1199.40,1121.76 1205.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,1110.00 C 1191.00,1121.76 1199.40,1121.76 1205.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,1110.00 C 1251.00,1121.76 1259.40,1121.76 1265.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,1110.00 C 1251.00,1121.76 1259.40,1121.76 1265.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,1110.00 C 1251.00,1121.76 1259.40,1121.76 1265.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,1110.00 C 1311.00,1121.76 1319.40,1121.76 1325.70,1110.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,1110.00 C 1311.00,1121.76 1319.40,1121.76 1325.70,1110.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,1110.00 C 1311.00,1121.76 1319.40,1121.76 1325.70,1110.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,1170.00 C 171.00,1181.76 179.40,1181.76 185.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,1170.00 C 171.00,1181.76 179.40,1181.76 185.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,1170.00 C 171.00,1181.76 179.40,1181.76 185.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,1170.00 C 231.00,1181.76 239.40,1181.76 245.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,1170.00 C 231.00,1181.76 239.40,1181.76 245.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,1170.00 C 231.00,1181.76 239.40,1181.76 245.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,1170.00 C 291.00,1181.76 299.40,1181.76 305.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,1170.00 C 291.00,1181.76 299.40,1181.76 305.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,1170.00 C 291.00,1181.76 299.40,1181.76 305.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,1170.00 C 351.00,1181.76 359.40,1181.76 365.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,1170.00 C 351.00,1181.76 359.40,1181.76 365.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,1170.00 C 351.00,1181.76 359.40,1181.76 365.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,1170.00 C 411.00,1181.76 419.40,1181.76 425.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,1170.00 C 411.00,1181.76 419.40,1181.76 425.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,1170.00 C 411.00,1181.76 419.40,1181.76 425.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,1170.00 C 471.00,1181.76 479.40,1181.76 485.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,1170.00 C 471.00,1181.76 479.40,1181.76 485.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,1170.00 C 471.00,1181.76 479.40,1181.76 485.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,1170.00 C 531.00,1181.76 539.40,1181.76 545.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,1170.00 C 531.00,1181.76 539.40,1181.76 545.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,1170.00 C 531.00,1181.76 539.40,1181.76 545.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,1170.00 C 591.00,1181.76 599.40,1181.76 605.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,1170.00 C 591.00,1181.76 599.40,1181.76 605.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,1170.00 C 591.00,1181.76 599.40,1181.76 605.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,1170.00 C 651.00,1181.76 659.40,1181.76 665.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,1170.00 C 651.00,1181.76 659.40,1181.76 665.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,1170.00 C 651.00,1181.76 659.40,1181.76 665.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,1170.00 C 711.00,1181.76 719.40,1181.76 725.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,1170.00 C 711.00,1181.76 719.40,1181.76 725.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,1170.00 C 711.00,1181.76 719.40,1181.76 725.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,1170.00 C 771.00,1181.76 779.40,1181.76 785.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,1170.00 C 771.00,1181.76 779.40,1181.76 785.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,1170.00 C 771.00,1181.76 779.40,1181.76 785.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,1170.00 C 831.00,1181.76 839.40,1181.76 845.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,1170.00 C 831.00,1181.76 839.40,1181.76 845.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,1170.00 C 831.00,1181.76 839.40,1181.76 845.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,1170.00 C 891.00,1181.76 899.40,1181.76 905.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,1170.00 C 891.00,1181.76 899.40,1181.76 905.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,1170.00 C 891.00,1181.76 899.40,1181.76 905.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,1170.00 C 951.00,1181.76 959.40,1181.76 965.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,1170.00 C 951.00,1181.76 959.40,1181.76 965.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,1170.00 C 951.00,1181.76 959.40,1181.76 965.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,1170.00 C 1011.00,1181.76 1019.40,1181.76 1025.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,1170.00 C 1011.00,1181.76 1019.40,1181.76 1025.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,1170.00 C 1011.00,1181.76 1019.40,1181.76 1025.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,1170.00 C 1071.00,1181.76 1079.40,1181.76 1085.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,1170.00 C 1071.00,1181.76 1079.40,1181.76 1085.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,1170.00 C 1071.00,1181.76 1079.40,1181.76 1085.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,1170.00 C 1131.00,1181.76 1139.40,1181.76 1145.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,1170.00 C 1131.00,1181.76 1139.40,1181.76 1145.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,1170.00 C 1131.00,1181.76 1139.40,1181.76 1145.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,1170.00 C 1191.00,1181.76 1199.40,1181.76 1205.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,1170.00 C 1191.00,1181.76 1199.40,1181.76 1205.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,1170.00 C 1191.00,1181.76 1199.40,1181.76 1205.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,1170.00 C 1251.00,1181.76 1259.40,1181.76 1265.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,1170.00 C 1251.00,1181.76 1259.40,1181.76 1265.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,1170.00 C 1251.00,1181.76 1259.40,1181.76 1265.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,1170.00 C 1311.00,1181.76 1319.40,1181.76 1325.70,1170.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,1170.00 C 1311.00,1181.76 1319.40,1181.76 1325.70,1170.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,1170.00 C 1311.00,1181.76 1319.40,1181.76 1325.70,1170.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,1230.00 C 171.00,1241.76 179.40,1241.76 185.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,1230.00 C 171.00,1241.76 179.40,1241.76 185.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,1230.00 C 171.00,1241.76 179.40,1241.76 185.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,1230.00 C 231.00,1241.76 239.40,1241.76 245.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,1230.00 C 231.00,1241.76 239.40,1241.76 245.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,1230.00 C 231.00,1241.76 239.40,1241.76 245.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,1230.00 C 291.00,1241.76 299.40,1241.76 305.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,1230.00 C 291.00,1241.76 299.40,1241.76 305.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,1230.00 C 291.00,1241.76 299.40,1241.76 305.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,1230.00 C 351.00,1241.76 359.40,1241.76 365.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,1230.00 C 351.00,1241.76 359.40,1241.76 365.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,1230.00 C 351.00,1241.76 359.40,1241.76 365.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,1230.00 C 411.00,1241.76 419.40,1241.76 425.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,1230.00 C 411.00,1241.76 419.40,1241.76 425.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,1230.00 C 411.00,1241.76 419.40,1241.76 425.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,1230.00 C 471.00,1241.76 479.40,1241.76 485.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,1230.00 C 471.00,1241.76 479.40,1241.76 485.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,1230.00 C 471.00,1241.76 479.40,1241.76 485.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,1230.00 C 531.00,1241.76 539.40,1241.76 545.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,1230.00 C 531.00,1241.76 539.40,1241.76 545.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,1230.00 C 531.00,1241.76 539.40,1241.76 545.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,1230.00 C 591.00,1241.76 599.40,1241.76 605.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,1230.00 C 591.00,1241.76 599.40,1241.76 605.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,1230.00 C 591.00,1241.76 599.40,1241.76 605.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,1230.00 C 651.00,1241.76 659.40,1241.76 665.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,1230.00 C 651.00,1241.76 659.40,1241.76 665.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,1230.00 C 651.00,1241.76 659.40,1241.76 665.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,1230.00 C 711.00,1241.76 719.40,1241.76 725.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,1230.00 C 711.00,1241.76 719.40,1241.76 725.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,1230.00 C 711.00,1241.76 719.40,1241.76 725.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,1230.00 C 771.00,1241.76 779.40,1241.76 785.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,1230.00 C 771.00,1241.76 779.40,1241.76 785.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,1230.00 C 771.00,1241.76 779.40,1241.76 785.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,1230.00 C 831.00,1241.76 839.40,1241.76 845.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,1230.00 C 831.00,1241.76 839.40,1241.76 845.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,1230.00 C 831.00,1241.76 839.40,1241.76 845.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,1230.00 C 891.00,1241.76 899.40,1241.76 905.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,1230.00 C 891.00,1241.76 899.40,1241.76 905.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,1230.00 C 891.00,1241.76 899.40,1241.76 905.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,1230.00 C 951.00,1241.76 959.40,1241.76 965.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,1230.00 C 951.00,1241.76 959.40,1241.76 965.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,1230.00 C 951.00,1241.76 959.40,1241.76 965.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,1230.00 C 1011.00,1241.76 1019.40,1241.76 1025.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,1230.00 C 1011.00,1241.76 1019.40,1241.76 1025.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,1230.00 C 1011.00,1241.76 1019.40,1241.76 1025.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,1230.00 C 1071.00,1241.76 1079.40,1241.76 1085.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,1230.00 C 1071.00,1241.76 1079.40,1241.76 1085.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,1230.00 C 1071.00,1241.76 1079.40,1241.76 1085.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,1230.00 C 1131.00,1241.76 1139.40,1241.76 1145.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,1230.00 C 1131.00,1241.76 1139.40,1241.76 1145.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,1230.00 C 1131.00,1241.76 1139.40,1241.76 1145.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,1230.00 C 1191.00,1241.76 1199.40,1241.76 1205.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,1230.00 C 1191.00,1241.76 1199.40,1241.76 1205.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,1230.00 C 1191.00,1241.76 1199.40,1241.76 1205.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,1230.00 C 1251.00,1241.76 1259.40,1241.76 1265.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,1230.00 C 1251.00,1241.76 1259.40,1241.76 1265.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,1230.00 C 1251.00,1241.76 1259.40,1241.76 1265.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,1230.00 C 1311.00,1241.76 1319.40,1241.76 1325.70,1230.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,1230.00 C 1311.00,1241.76 1319.40,1241.76 1325.70,1230.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,1230.00 C 1311.00,1241.76 1319.40,1241.76 1325.70,1230.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,1290.00 C 171.00,1301.76 179.40,1301.76 185.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,1290.00 C 171.00,1301.76 179.40,1301.76 185.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,1290.00 C 171.00,1301.76 179.40,1301.76 185.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,1290.00 C 231.00,1301.76 239.40,1301.76 245.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,1290.00 C 231.00,1301.76 239.40,1301.76 245.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,1290.00 C 231.00,1301.76 239.40,1301.76 245.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,1290.00 C 291.00,1301.76 299.40,1301.76 305.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,1290.00 C 291.00,1301.76 299.40,1301.76 305.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,1290.00 C 291.00,1301.76 299.40,1301.76 305.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,1290.00 C 351.00,1301.76 359.40,1301.76 365.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,1290.00 C 351.00,1301.76 359.40,1301.76 365.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,1290.00 C 351.00,1301.76 359.40,1301.76 365.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,1290.00 C 411.00,1301.76 419.40,1301.76 425.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,1290.00 C 411.00,1301.76 419.40,1301.76 425.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,1290.00 C 411.00,1301.76 419.40,1301.76 425.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,1290.00 C 471.00,1301.76 479.40,1301.76 485.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,1290.00 C 471.00,1301.76 479.40,1301.76 485.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,1290.00 C 471.00,1301.76 479.40,1301.76 485.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,1290.00 C 531.00,1301.76 539.40,1301.76 545.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,1290.00 C 531.00,1301.76 539.40,1301.76 545.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,1290.00 C 531.00,1301.76 539.40,1301.76 545.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,1290.00 C 591.00,1301.76 599.40,1301.76 605.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,1290.00 C 591.00,1301.76 599.40,1301.76 605.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,1290.00 C 591.00,1301.76 599.40,1301.76 605.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,1290.00 C 651.00,1301.76 659.40,1301.76 665.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,1290.00 C 651.00,1301.76 659.40,1301.76 665.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,1290.00 C 651.00,1301.76 659.40,1301.76 665.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,1290.00 C 711.00,1301.76 719.40,1301.76 725.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,1290.00 C 711.00,1301.76 719.40,1301.76 725.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,1290.00 C 711.00,1301.76 719.40,1301.76 725.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,1290.00 C 771.00,1301.76 779.40,1301.76 785.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,1290.00 C 771.00,1301.76 779.40,1301.76 785.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,1290.00 C 771.00,1301.76 779.40,1301.76 785.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,1290.00 C 831.00,1301.76 839.40,1301.76 845.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,1290.00 C 831.00,1301.76 839.40,1301.76 845.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,1290.00 C 831.00,1301.76 839.40,1301.76 845.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,1290.00 C 891.00,1301.76 899.40,1301.76 905.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,1290.00 C 891.00,1301.76 899.40,1301.76 905.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,1290.00 C 891.00,1301.76 899.40,1301.76 905.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,1290.00 C 951.00,1301.76 959.40,1301.76 965.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,1290.00 C 951.00,1301.76 959.40,1301.76 965.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,1290.00 C 951.00,1301.76 959.40,1301.76 965.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,1290.00 C 1011.00,1301.76 1019.40,1301.76 1025.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,1290.00 C 1011.00,1301.76 1019.40,1301.76 1025.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,1290.00 C 1011.00,1301.76 1019.40,1301.76 1025.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,1290.00 C 1071.00,1301.76 1079.40,1301.76 1085.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,1290.00 C 1071.00,1301.76 1079.40,1301.76 1085.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,1290.00 C 1071.00,1301.76 1079.40,1301.76 1085.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,1290.00 C 1131.00,1301.76 1139.40,1301.76 1145.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,1290.00 C 1131.00,1301.76 1139.40,1301.76 1145.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,1290.00 C 1131.00,1301.76 1139.40,1301.76 1145.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,1290.00 C 1191.00,1301.76 1199.40,1301.76 1205.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,1290.00 C 1191.00,1301.76 1199.40,1301.76 1205.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,1290.00 C 1191.00,1301.76 1199.40,1301.76 1205.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,1290.00 C 1251.00,1301.76 1259.40,1301.76 1265.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,1290.00 C 1251.00,1301.76 1259.40,1301.76 1265.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,1290.00 C 1251.00,1301.76 1259.40,1301.76 1265.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,1290.00 C 1311.00,1301.76 1319.40,1301.76 1325.70,1290.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,1290.00 C 1311.00,1301.76 1319.40,1301.76 1325.70,1290.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,1290.00 C 1311.00,1301.76 1319.40,1301.76 1325.70,1290.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 164.70,1350.00 C 171.00,1361.76 179.40,1361.76 185.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 164.70,1350.00 C 171.00,1361.76 179.40,1361.76 185.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 164.70,1350.00 C 171.00,1361.76 179.40,1361.76 185.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 224.70,1350.00 C 231.00,1361.76 239.40,1361.76 245.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 224.70,1350.00 C 231.00,1361.76 239.40,1361.76 245.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 224.70,1350.00 C 231.00,1361.76 239.40,1361.76 245.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 284.70,1350.00 C 291.00,1361.76 299.40,1361.76 305.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 284.70,1350.00 C 291.00,1361.76 299.40,1361.76 305.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 284.70,1350.00 C 291.00,1361.76 299.40,1361.76 305.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 344.70,1350.00 C 351.00,1361.76 359.40,1361.76 365.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 344.70,1350.00 C 351.00,1361.76 359.40,1361.76 365.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 344.70,1350.00 C 351.00,1361.76 359.40,1361.76 365.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 404.70,1350.00 C 411.00,1361.76 419.40,1361.76 425.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 404.70,1350.00 C 411.00,1361.76 419.40,1361.76 425.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 404.70,1350.00 C 411.00,1361.76 419.40,1361.76 425.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 464.70,1350.00 C 471.00,1361.76 479.40,1361.76 485.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 464.70,1350.00 C 471.00,1361.76 479.40,1361.76 485.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 464.70,1350.00 C 471.00,1361.76 479.40,1361.76 485.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 524.70,1350.00 C 531.00,1361.76 539.40,1361.76 545.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 524.70,1350.00 C 531.00,1361.76 539.40,1361.76 545.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 524.70,1350.00 C 531.00,1361.76 539.40,1361.76 545.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 584.70,1350.00 C 591.00,1361.76 599.40,1361.76 605.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 584.70,1350.00 C 591.00,1361.76 599.40,1361.76 605.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 584.70,1350.00 C 591.00,1361.76 599.40,1361.76 605.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 644.70,1350.00 C 651.00,1361.76 659.40,1361.76 665.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 644.70,1350.00 C 651.00,1361.76 659.40,1361.76 665.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 644.70,1350.00 C 651.00,1361.76 659.40,1361.76 665.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 704.70,1350.00 C 711.00,1361.76 719.40,1361.76 725.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 704.70,1350.00 C 711.00,1361.76 719.40,1361.76 725.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 704.70,1350.00 C 711.00,1361.76 719.40,1361.76 725.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 764.70,1350.00 C 771.00,1361.76 779.40,1361.76 785.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 764.70,1350.00 C 771.00,1361.76 779.40,1361.76 785.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 764.70,1350.00 C 771.00,1361.76 779.40,1361.76 785.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 824.70,1350.00 C 831.00,1361.76 839.40,1361.76 845.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 824.70,1350.00 C 831.00,1361.76 839.40,1361.76 845.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 824.70,1350.00 C 831.00,1361.76 839.40,1361.76 845.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 884.70,1350.00 C 891.00,1361.76 899.40,1361.76 905.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 884.70,1350.00 C 891.00,1361.76 899.40,1361.76 905.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 884.70,1350.00 C 891.00,1361.76 899.40,1361.76 905.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 944.70,1350.00 C 951.00,1361.76 959.40,1361.76 965.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 944.70,1350.00 C 951.00,1361.76 959.40,1361.76 965.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 944.70,1350.00 C 951.00,1361.76 959.40,1361.76 965.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1004.70,1350.00 C 1011.00,1361.76 1019.40,1361.76 1025.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1004.70,1350.00 C 1011.00,1361.76 1019.40,1361.76 1025.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1004.70,1350.00 C 1011.00,1361.76 1019.40,1361.76 1025.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1064.70,1350.00 C 1071.00,1361.76 1079.40,1361.76 1085.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1064.70,1350.00 C 1071.00,1361.76 1079.40,1361.76 1085.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1064.70,1350.00 C 1071.00,1361.76 1079.40,1361.76 1085.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1124.70,1350.00 C 1131.00,1361.76 1139.40,1361.76 1145.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1124.70,1350.00 C 1131.00,1361.76 1139.40,1361.76 1145.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1124.70,1350.00 C 1131.00,1361.76 1139.40,1361.76 1145.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1184.70,1350.00 C 1191.00,1361.76 1199.40,1361.76 1205.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1184.70,1350.00 C 1191.00,1361.76 1199.40,1361.76 1205.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1184.70,1350.00 C 1191.00,1361.76 1199.40,1361.76 1205.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1244.70,1350.00 C 1251.00,1361.76 1259.40,1361.76 1265.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1244.70,1350.00 C 1251.00,1361.76 1259.40,1361.76 1265.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1244.70,1350.00 C 1251.00,1361.76 1259.40,1361.76 1265.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1304.70,1350.00 C 1311.00,1361.76 1319.40,1361.76 1325.70,1350.00" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1304.70,1350.00 C 1311.00,1361.76 1319.40,1361.76 1325.70,1350.00" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1304.70,1350.00 C 1311.00,1361.76 1319.40,1361.76 1325.70,1350.00" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,164.70 C 138.24,171.00 138.24,179.40 150.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,164.70 C 138.24,171.00 138.24,179.40 150.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,164.70 C 138.24,171.00 138.24,179.40 150.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,164.70 C 198.24,171.00 198.24,179.40 210.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,164.70 C 198.24,171.00 198.24,179.40 210.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,164.70 C 198.24,171.00 198.24,179.40 210.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,164.70 C 258.24,171.00 258.24,179.40 270.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,164.70 C 258.24,171.00 258.24,179.40 270.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,164.70 C 258.24,171.00 258.24,179.40 270.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,164.70 C 318.24,171.00 318.24,179.40 330.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,164.70 C 318.24,171.00 318.24,179.40 330.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,164.70 C 318.24,171.00 318.24,179.40 330.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,164.70 C 378.24,171.00 378.24,179.40 390.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,164.70 C 378.24,171.00 378.24,179.40 390.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,164.70 C 378.24,171.00 378.24,179.40 390.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,164.70 C 438.24,171.00 438.24,179.40 450.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,164.70 C 438.24,171.00 438.24,179.40 450.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,164.70 C 438.24,171.00 438.24,179.40 450.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,164.70 C 498.24,171.00 498.24,179.40 510.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,164.70 C 498.24,171.00 498.24,179.40 510.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,164.70 C 498.24,171.00 498.24,179.40 510.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,164.70 C 558.24,171.00 558.24,179.40 570.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,164.70 C 558.24,171.00 558.24,179.40 570.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,164.70 C 558.24,171.00 558.24,179.40 570.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,164.70 C 618.24,171.00 618.24,179.40 630.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,164.70 C 618.24,171.00 618.24,179.40 630.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,164.70 C 618.24,171.00 618.24,179.40 630.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,164.70 C 678.24,171.00 678.24,179.40 690.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,164.70 C 678.24,171.00 678.24,179.40 690.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,164.70 C 678.24,171.00 678.24,179.40 690.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,164.70 C 738.24,171.00 738.24,179.40 750.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,164.70 C 738.24,171.00 738.24,179.40 750.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,164.70 C 738.24,171.00 738.24,179.40 750.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,164.70 C 798.24,171.00 798.24,179.40 810.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,164.70 C 798.24,171.00 798.24,179.40 810.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,164.70 C 798.24,171.00 798.24,179.40 810.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,164.70 C 858.24,171.00 858.24,179.40 870.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,164.70 C 858.24,171.00 858.24,179.40 870.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,164.70 C 858.24,171.00 858.24,179.40 870.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,164.70 C 918.24,171.00 918.24,179.40 930.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,164.70 C 918.24,171.00 918.24,179.40 930.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,164.70 C 918.24,171.00 918.24,179.40 930.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,164.70 C 978.24,171.00 978.24,179.40 990.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,164.70 C 978.24,171.00 978.24,179.40 990.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,164.70 C 978.24,171.00 978.24,179.40 990.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,164.70 C 1038.24,171.00 1038.24,179.40 1050.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,164.70 C 1038.24,171.00 1038.24,179.40 1050.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,164.70 C 1038.24,171.00 1038.24,179.40 1050.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,164.70 C 1098.24,171.00 1098.24,179.40 1110.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,164.70 C 1098.24,171.00 1098.24,179.40 1110.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,164.70 C 1098.24,171.00 1098.24,179.40 1110.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,164.70 C 1158.24,171.00 1158.24,179.40 1170.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,164.70 C 1158.24,171.00 1158.24,179.40 1170.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,164.70 C 1158.24,171.00 1158.24,179.40 1170.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,164.70 C 1218.24,171.00 1218.24,179.40 1230.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,164.70 C 1218.24,171.00 1218.24,179.40 1230.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,164.70 C 1218.24,171.00 1218.24,179.40 1230.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,164.70 C 1278.24,171.00 1278.24,179.40 1290.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,164.70 C 1278.24,171.00 1278.24,179.40 1290.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,164.70 C 1278.24,171.00 1278.24,179.40 1290.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,164.70 C 1338.24,171.00 1338.24,179.40 1350.00,185.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,164.70 C 1338.24,171.00 1338.24,179.40 1350.00,185.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,164.70 C 1338.24,171.00 1338.24,179.40 1350.00,185.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,224.70 C 138.24,231.00 138.24,239.40 150.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,224.70 C 138.24,231.00 138.24,239.40 150.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,224.70 C 138.24,231.00 138.24,239.40 150.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,224.70 C 198.24,231.00 198.24,239.40 210.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,224.70 C 198.24,231.00 198.24,239.40 210.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,224.70 C 198.24,231.00 198.24,239.40 210.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,224.70 C 258.24,231.00 258.24,239.40 270.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,224.70 C 258.24,231.00 258.24,239.40 270.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,224.70 C 258.24,231.00 258.24,239.40 270.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,224.70 C 318.24,231.00 318.24,239.40 330.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,224.70 C 318.24,231.00 318.24,239.40 330.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,224.70 C 318.24,231.00 318.24,239.40 330.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,224.70 C 378.24,231.00 378.24,239.40 390.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,224.70 C 378.24,231.00 378.24,239.40 390.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,224.70 C 378.24,231.00 378.24,239.40 390.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,224.70 C 438.24,231.00 438.24,239.40 450.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,224.70 C 438.24,231.00 438.24,239.40 450.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,224.70 C 438.24,231.00 438.24,239.40 450.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,224.70 C 498.24,231.00 498.24,239.40 510.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,224.70 C 498.24,231.00 498.24,239.40 510.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,224.70 C 498.24,231.00 498.24,239.40 510.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,224.70 C 558.24,231.00 558.24,239.40 570.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,224.70 C 558.24,231.00 558.24,239.40 570.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,224.70 C 558.24,231.00 558.24,239.40 570.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,224.70 C 618.24,231.00 618.24,239.40 630.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,224.70 C 618.24,231.00 618.24,239.40 630.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,224.70 C 618.24,231.00 618.24,239.40 630.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,224.70 C 678.24,231.00 678.24,239.40 690.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,224.70 C 678.24,231.00 678.24,239.40 690.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,224.70 C 678.24,231.00 678.24,239.40 690.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,224.70 C 738.24,231.00 738.24,239.40 750.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,224.70 C 738.24,231.00 738.24,239.40 750.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,224.70 C 738.24,231.00 738.24,239.40 750.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,224.70 C 798.24,231.00 798.24,239.40 810.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,224.70 C 798.24,231.00 798.24,239.40 810.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,224.70 C 798.24,231.00 798.24,239.40 810.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,224.70 C 858.24,231.00 858.24,239.40 870.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,224.70 C 858.24,231.00 858.24,239.40 870.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,224.70 C 858.24,231.00 858.24,239.40 870.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,224.70 C 918.24,231.00 918.24,239.40 930.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,224.70 C 918.24,231.00 918.24,239.40 930.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,224.70 C 918.24,231.00 918.24,239.40 930.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,224.70 C 978.24,231.00 978.24,239.40 990.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,224.70 C 978.24,231.00 978.24,239.40 990.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,224.70 C 978.24,231.00 978.24,239.40 990.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,224.70 C 1038.24,231.00 1038.24,239.40 1050.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,224.70 C 1038.24,231.00 1038.24,239.40 1050.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,224.70 C 1038.24,231.00 1038.24,239.40 1050.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,224.70 C 1098.24,231.00 1098.24,239.40 1110.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,224.70 C 1098.24,231.00 1098.24,239.40 1110.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,224.70 C 1098.24,231.00 1098.24,239.40 1110.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,224.70 C 1158.24,231.00 1158.24,239.40 1170.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,224.70 C 1158.24,231.00 1158.24,239.40 1170.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,224.70 C 1158.24,231.00 1158.24,239.40 1170.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,224.70 C 1218.24,231.00 1218.24,239.40 1230.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,224.70 C 1218.24,231.00 1218.24,239.40 1230.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,224.70 C 1218.24,231.00 1218.24,239.40 1230.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,224.70 C 1278.24,231.00 1278.24,239.40 1290.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,224.70 C 1278.24,231.00 1278.24,239.40 1290.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,224.70 C 1278.24,231.00 1278.24,239.40 1290.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,224.70 C 1338.24,231.00 1338.24,239.40 1350.00,245.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,224.70 C 1338.24,231.00 1338.24,239.40 1350.00,245.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,224.70 C 1338.24,231.00 1338.24,239.40 1350.00,245.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,284.70 C 138.24,291.00 138.24,299.40 150.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,284.70 C 138.24,291.00 138.24,299.40 150.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,284.70 C 138.24,291.00 138.24,299.40 150.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,284.70 C 198.24,291.00 198.24,299.40 210.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,284.70 C 198.24,291.00 198.24,299.40 210.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,284.70 C 198.24,291.00 198.24,299.40 210.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,284.70 C 258.24,291.00 258.24,299.40 270.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,284.70 C 258.24,291.00 258.24,299.40 270.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,284.70 C 258.24,291.00 258.24,299.40 270.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,284.70 C 318.24,291.00 318.24,299.40 330.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,284.70 C 318.24,291.00 318.24,299.40 330.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,284.70 C 318.24,291.00 318.24,299.40 330.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,284.70 C 378.24,291.00 378.24,299.40 390.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,284.70 C 378.24,291.00 378.24,299.40 390.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,284.70 C 378.24,291.00 378.24,299.40 390.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,284.70 C 438.24,291.00 438.24,299.40 450.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,284.70 C 438.24,291.00 438.24,299.40 450.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,284.70 C 438.24,291.00 438.24,299.40 450.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,284.70 C 498.24,291.00 498.24,299.40 510.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,284.70 C 498.24,291.00 498.24,299.40 510.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,284.70 C 498.24,291.00 498.24,299.40 510.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,284.70 C 558.24,291.00 558.24,299.40 570.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,284.70 C 558.24,291.00 558.24,299.40 570.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,284.70 C 558.24,291.00 558.24,299.40 570.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,284.70 C 618.24,291.00 618.24,299.40 630.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,284.70 C 618.24,291.00 618.24,299.40 630.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,284.70 C 618.24,291.00 618.24,299.40 630.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,284.70 C 678.24,291.00 678.24,299.40 690.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,284.70 C 678.24,291.00 678.24,299.40 690.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,284.70 C 678.24,291.00 678.24,299.40 690.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,284.70 C 738.24,291.00 738.24,299.40 750.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,284.70 C 738.24,291.00 738.24,299.40 750.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,284.70 C 738.24,291.00 738.24,299.40 750.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,284.70 C 798.24,291.00 798.24,299.40 810.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,284.70 C 798.24,291.00 798.24,299.40 810.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,284.70 C 798.24,291.00 798.24,299.40 810.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,284.70 C 858.24,291.00 858.24,299.40 870.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,284.70 C 858.24,291.00 858.24,299.40 870.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,284.70 C 858.24,291.00 858.24,299.40 870.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,284.70 C 918.24,291.00 918.24,299.40 930.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,284.70 C 918.24,291.00 918.24,299.40 930.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,284.70 C 918.24,291.00 918.24,299.40 930.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,284.70 C 978.24,291.00 978.24,299.40 990.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,284.70 C 978.24,291.00 978.24,299.40 990.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,284.70 C 978.24,291.00 978.24,299.40 990.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,284.70 C 1038.24,291.00 1038.24,299.40 1050.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,284.70 C 1038.24,291.00 1038.24,299.40 1050.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,284.70 C 1038.24,291.00 1038.24,299.40 1050.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,284.70 C 1098.24,291.00 1098.24,299.40 1110.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,284.70 C 1098.24,291.00 1098.24,299.40 1110.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,284.70 C 1098.24,291.00 1098.24,299.40 1110.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,284.70 C 1158.24,291.00 1158.24,299.40 1170.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,284.70 C 1158.24,291.00 1158.24,299.40 1170.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,284.70 C 1158.24,291.00 1158.24,299.40 1170.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,284.70 C 1218.24,291.00 1218.24,299.40 1230.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,284.70 C 1218.24,291.00 1218.24,299.40 1230.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,284.70 C 1218.24,291.00 1218.24,299.40 1230.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,284.70 C 1278.24,291.00 1278.24,299.40 1290.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,284.70 C 1278.24,291.00 1278.24,299.40 1290.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,284.70 C 1278.24,291.00 1278.24,299.40 1290.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,284.70 C 1338.24,291.00 1338.24,299.40 1350.00,305.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,284.70 C 1338.24,291.00 1338.24,299.40 1350.00,305.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,284.70 C 1338.24,291.00 1338.24,299.40 1350.00,305.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,344.70 C 138.24,351.00 138.24,359.40 150.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,344.70 C 138.24,351.00 138.24,359.40 150.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,344.70 C 138.24,351.00 138.24,359.40 150.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,344.70 C 198.24,351.00 198.24,359.40 210.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,344.70 C 198.24,351.00 198.24,359.40 210.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,344.70 C 198.24,351.00 198.24,359.40 210.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,344.70 C 258.24,351.00 258.24,359.40 270.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,344.70 C 258.24,351.00 258.24,359.40 270.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,344.70 C 258.24,351.00 258.24,359.40 270.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,344.70 C 318.24,351.00 318.24,359.40 330.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,344.70 C 318.24,351.00 318.24,359.40 330.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,344.70 C 318.24,351.00 318.24,359.40 330.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,344.70 C 378.24,351.00 378.24,359.40 390.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,344.70 C 378.24,351.00 378.24,359.40 390.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,344.70 C 378.24,351.00 378.24,359.40 390.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,344.70 C 438.24,351.00 438.24,359.40 450.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,344.70 C 438.24,351.00 438.24,359.40 450.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,344.70 C 438.24,351.00 438.24,359.40 450.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,344.70 C 498.24,351.00 498.24,359.40 510.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,344.70 C 498.24,351.00 498.24,359.40 510.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,344.70 C 498.24,351.00 498.24,359.40 510.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,344.70 C 558.24,351.00 558.24,359.40 570.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,344.70 C 558.24,351.00 558.24,359.40 570.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,344.70 C 558.24,351.00 558.24,359.40 570.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,344.70 C 618.24,351.00 618.24,359.40 630.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,344.70 C 618.24,351.00 618.24,359.40 630.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,344.70 C 618.24,351.00 618.24,359.40 630.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,344.70 C 678.24,351.00 678.24,359.40 690.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,344.70 C 678.24,351.00 678.24,359.40 690.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,344.70 C 678.24,351.00 678.24,359.40 690.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,344.70 C 738.24,351.00 738.24,359.40 750.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,344.70 C 738.24,351.00 738.24,359.40 750.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,344.70 C 738.24,351.00 738.24,359.40 750.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,344.70 C 798.24,351.00 798.24,359.40 810.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,344.70 C 798.24,351.00 798.24,359.40 810.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,344.70 C 798.24,351.00 798.24,359.40 810.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,344.70 C 858.24,351.00 858.24,359.40 870.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,344.70 C 858.24,351.00 858.24,359.40 870.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,344.70 C 858.24,351.00 858.24,359.40 870.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,344.70 C 918.24,351.00 918.24,359.40 930.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,344.70 C 918.24,351.00 918.24,359.40 930.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,344.70 C 918.24,351.00 918.24,359.40 930.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,344.70 C 978.24,351.00 978.24,359.40 990.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,344.70 C 978.24,351.00 978.24,359.40 990.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,344.70 C 978.24,351.00 978.24,359.40 990.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,344.70 C 1038.24,351.00 1038.24,359.40 1050.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,344.70 C 1038.24,351.00 1038.24,359.40 1050.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,344.70 C 1038.24,351.00 1038.24,359.40 1050.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,344.70 C 1098.24,351.00 1098.24,359.40 1110.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,344.70 C 1098.24,351.00 1098.24,359.40 1110.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,344.70 C 1098.24,351.00 1098.24,359.40 1110.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,344.70 C 1158.24,351.00 1158.24,359.40 1170.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,344.70 C 1158.24,351.00 1158.24,359.40 1170.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,344.70 C 1158.24,351.00 1158.24,359.40 1170.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,344.70 C 1218.24,351.00 1218.24,359.40 1230.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,344.70 C 1218.24,351.00 1218.24,359.40 1230.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,344.70 C 1218.24,351.00 1218.24,359.40 1230.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,344.70 C 1278.24,351.00 1278.24,359.40 1290.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,344.70 C 1278.24,351.00 1278.24,359.40 1290.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,344.70 C 1278.24,351.00 1278.24,359.40 1290.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,344.70 C 1338.24,351.00 1338.24,359.40 1350.00,365.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,344.70 C 1338.24,351.00 1338.24,359.40 1350.00,365.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,344.70 C 1338.24,351.00 1338.24,359.40 1350.00,365.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,404.70 C 138.24,411.00 138.24,419.40 150.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,404.70 C 138.24,411.00 138.24,419.40 150.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,404.70 C 138.24,411.00 138.24,419.40 150.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,404.70 C 198.24,411.00 198.24,419.40 210.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,404.70 C 198.24,411.00 198.24,419.40 210.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,404.70 C 198.24,411.00 198.24,419.40 210.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,404.70 C 258.24,411.00 258.24,419.40 270.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,404.70 C 258.24,411.00 258.24,419.40 270.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,404.70 C 258.24,411.00 258.24,419.40 270.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,404.70 C 318.24,411.00 318.24,419.40 330.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,404.70 C 318.24,411.00 318.24,419.40 330.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,404.70 C 318.24,411.00 318.24,419.40 330.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,404.70 C 378.24,411.00 378.24,419.40 390.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,404.70 C 378.24,411.00 378.24,419.40 390.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,404.70 C 378.24,411.00 378.24,419.40 390.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,404.70 C 438.24,411.00 438.24,419.40 450.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,404.70 C 438.24,411.00 438.24,419.40 450.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,404.70 C 438.24,411.00 438.24,419.40 450.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,404.70 C 498.24,411.00 498.24,419.40 510.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,404.70 C 498.24,411.00 498.24,419.40 510.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,404.70 C 498.24,411.00 498.24,419.40 510.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,404.70 C 558.24,411.00 558.24,419.40 570.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,404.70 C 558.24,411.00 558.24,419.40 570.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,404.70 C 558.24,411.00 558.24,419.40 570.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,404.70 C 618.24,411.00 618.24,419.40 630.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,404.70 C 618.24,411.00 618.24,419.40 630.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,404.70 C 618.24,411.00 618.24,419.40 630.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,404.70 C 678.24,411.00 678.24,419.40 690.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,404.70 C 678.24,411.00 678.24,419.40 690.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,404.70 C 678.24,411.00 678.24,419.40 690.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,404.70 C 738.24,411.00 738.24,419.40 750.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,404.70 C 738.24,411.00 738.24,419.40 750.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,404.70 C 738.24,411.00 738.24,419.40 750.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,404.70 C 798.24,411.00 798.24,419.40 810.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,404.70 C 798.24,411.00 798.24,419.40 810.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,404.70 C 798.24,411.00 798.24,419.40 810.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,404.70 C 858.24,411.00 858.24,419.40 870.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,404.70 C 858.24,411.00 858.24,419.40 870.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,404.70 C 858.24,411.00 858.24,419.40 870.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,404.70 C 918.24,411.00 918.24,419.40 930.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,404.70 C 918.24,411.00 918.24,419.40 930.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,404.70 C 918.24,411.00 918.24,419.40 930.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,404.70 C 978.24,411.00 978.24,419.40 990.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,404.70 C 978.24,411.00 978.24,419.40 990.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,404.70 C 978.24,411.00 978.24,419.40 990.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,404.70 C 1038.24,411.00 1038.24,419.40 1050.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,404.70 C 1038.24,411.00 1038.24,419.40 1050.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,404.70 C 1038.24,411.00 1038.24,419.40 1050.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,404.70 C 1098.24,411.00 1098.24,419.40 1110.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,404.70 C 1098.24,411.00 1098.24,419.40 1110.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,404.70 C 1098.24,411.00 1098.24,419.40 1110.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,404.70 C 1158.24,411.00 1158.24,419.40 1170.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,404.70 C 1158.24,411.00 1158.24,419.40 1170.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,404.70 C 1158.24,411.00 1158.24,419.40 1170.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,404.70 C 1218.24,411.00 1218.24,419.40 1230.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,404.70 C 1218.24,411.00 1218.24,419.40 1230.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,404.70 C 1218.24,411.00 1218.24,419.40 1230.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,404.70 C 1278.24,411.00 1278.24,419.40 1290.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,404.70 C 1278.24,411.00 1278.24,419.40 1290.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,404.70 C 1278.24,411.00 1278.24,419.40 1290.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,404.70 C 1338.24,411.00 1338.24,419.40 1350.00,425.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,404.70 C 1338.24,411.00 1338.24,419.40 1350.00,425.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,404.70 C 1338.24,411.00 1338.24,419.40 1350.00,425.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,464.70 C 138.24,471.00 138.24,479.40 150.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,464.70 C 138.24,471.00 138.24,479.40 150.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,464.70 C 138.24,471.00 138.24,479.40 150.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,464.70 C 198.24,471.00 198.24,479.40 210.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,464.70 C 198.24,471.00 198.24,479.40 210.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,464.70 C 198.24,471.00 198.24,479.40 210.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,464.70 C 258.24,471.00 258.24,479.40 270.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,464.70 C 258.24,471.00 258.24,479.40 270.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,464.70 C 258.24,471.00 258.24,479.40 270.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,464.70 C 318.24,471.00 318.24,479.40 330.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,464.70 C 318.24,471.00 318.24,479.40 330.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,464.70 C 318.24,471.00 318.24,479.40 330.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,464.70 C 378.24,471.00 378.24,479.40 390.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,464.70 C 378.24,471.00 378.24,479.40 390.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,464.70 C 378.24,471.00 378.24,479.40 390.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,464.70 C 438.24,471.00 438.24,479.40 450.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,464.70 C 438.24,471.00 438.24,479.40 450.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,464.70 C 438.24,471.00 438.24,479.40 450.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,464.70 C 498.24,471.00 498.24,479.40 510.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,464.70 C 498.24,471.00 498.24,479.40 510.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,464.70 C 498.24,471.00 498.24,479.40 510.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,464.70 C 558.24,471.00 558.24,479.40 570.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,464.70 C 558.24,471.00 558.24,479.40 570.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,464.70 C 558.24,471.00 558.24,479.40 570.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,464.70 C 618.24,471.00 618.24,479.40 630.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,464.70 C 618.24,471.00 618.24,479.40 630.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,464.70 C 618.24,471.00 618.24,479.40 630.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,464.70 C 678.24,471.00 678.24,479.40 690.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,464.70 C 678.24,471.00 678.24,479.40 690.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,464.70 C 678.24,471.00 678.24,479.40 690.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,464.70 C 738.24,471.00 738.24,479.40 750.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,464.70 C 738.24,471.00 738.24,479.40 750.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,464.70 C 738.24,471.00 738.24,479.40 750.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,464.70 C 798.24,471.00 798.24,479.40 810.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,464.70 C 798.24,471.00 798.24,479.40 810.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,464.70 C 798.24,471.00 798.24,479.40 810.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,464.70 C 858.24,471.00 858.24,479.40 870.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,464.70 C 858.24,471.00 858.24,479.40 870.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,464.70 C 858.24,471.00 858.24,479.40 870.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,464.70 C 918.24,471.00 918.24,479.40 930.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,464.70 C 918.24,471.00 918.24,479.40 930.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,464.70 C 918.24,471.00 918.24,479.40 930.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,464.70 C 978.24,471.00 978.24,479.40 990.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,464.70 C 978.24,471.00 978.24,479.40 990.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,464.70 C 978.24,471.00 978.24,479.40 990.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,464.70 C 1038.24,471.00 1038.24,479.40 1050.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,464.70 C 1038.24,471.00 1038.24,479.40 1050.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,464.70 C 1038.24,471.00 1038.24,479.40 1050.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,464.70 C 1098.24,471.00 1098.24,479.40 1110.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,464.70 C 1098.24,471.00 1098.24,479.40 1110.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,464.70 C 1098.24,471.00 1098.24,479.40 1110.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,464.70 C 1158.24,471.00 1158.24,479.40 1170.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,464.70 C 1158.24,471.00 1158.24,479.40 1170.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,464.70 C 1158.24,471.00 1158.24,479.40 1170.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,464.70 C 1218.24,471.00 1218.24,479.40 1230.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,464.70 C 1218.24,471.00 1218.24,479.40 1230.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,464.70 C 1218.24,471.00 1218.24,479.40 1230.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,464.70 C 1278.24,471.00 1278.24,479.40 1290.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,464.70 C 1278.24,471.00 1278.24,479.40 1290.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,464.70 C 1278.24,471.00 1278.24,479.40 1290.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,464.70 C 1338.24,471.00 1338.24,479.40 1350.00,485.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,464.70 C 1338.24,471.00 1338.24,479.40 1350.00,485.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,464.70 C 1338.24,471.00 1338.24,479.40 1350.00,485.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,524.70 C 138.24,531.00 138.24,539.40 150.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,524.70 C 138.24,531.00 138.24,539.40 150.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,524.70 C 138.24,531.00 138.24,539.40 150.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,524.70 C 198.24,531.00 198.24,539.40 210.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,524.70 C 198.24,531.00 198.24,539.40 210.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,524.70 C 198.24,531.00 198.24,539.40 210.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,524.70 C 258.24,531.00 258.24,539.40 270.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,524.70 C 258.24,531.00 258.24,539.40 270.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,524.70 C 258.24,531.00 258.24,539.40 270.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,524.70 C 318.24,531.00 318.24,539.40 330.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,524.70 C 318.24,531.00 318.24,539.40 330.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,524.70 C 318.24,531.00 318.24,539.40 330.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,524.70 C 378.24,531.00 378.24,539.40 390.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,524.70 C 378.24,531.00 378.24,539.40 390.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,524.70 C 378.24,531.00 378.24,539.40 390.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,524.70 C 438.24,531.00 438.24,539.40 450.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,524.70 C 438.24,531.00 438.24,539.40 450.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,524.70 C 438.24,531.00 438.24,539.40 450.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,524.70 C 498.24,531.00 498.24,539.40 510.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,524.70 C 498.24,531.00 498.24,539.40 510.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,524.70 C 498.24,531.00 498.24,539.40 510.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,524.70 C 558.24,531.00 558.24,539.40 570.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,524.70 C 558.24,531.00 558.24,539.40 570.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,524.70 C 558.24,531.00 558.24,539.40 570.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,524.70 C 618.24,531.00 618.24,539.40 630.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,524.70 C 618.24,531.00 618.24,539.40 630.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,524.70 C 618.24,531.00 618.24,539.40 630.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,524.70 C 678.24,531.00 678.24,539.40 690.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,524.70 C 678.24,531.00 678.24,539.40 690.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,524.70 C 678.24,531.00 678.24,539.40 690.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,524.70 C 738.24,531.00 738.24,539.40 750.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,524.70 C 738.24,531.00 738.24,539.40 750.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,524.70 C 738.24,531.00 738.24,539.40 750.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,524.70 C 798.24,531.00 798.24,539.40 810.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,524.70 C 798.24,531.00 798.24,539.40 810.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,524.70 C 798.24,531.00 798.24,539.40 810.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,524.70 C 858.24,531.00 858.24,539.40 870.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,524.70 C 858.24,531.00 858.24,539.40 870.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,524.70 C 858.24,531.00 858.24,539.40 870.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,524.70 C 918.24,531.00 918.24,539.40 930.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,524.70 C 918.24,531.00 918.24,539.40 930.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,524.70 C 918.24,531.00 918.24,539.40 930.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,524.70 C 978.24,531.00 978.24,539.40 990.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,524.70 C 978.24,531.00 978.24,539.40 990.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,524.70 C 978.24,531.00 978.24,539.40 990.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,524.70 C 1038.24,531.00 1038.24,539.40 1050.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,524.70 C 1038.24,531.00 1038.24,539.40 1050.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,524.70 C 1038.24,531.00 1038.24,539.40 1050.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,524.70 C 1098.24,531.00 1098.24,539.40 1110.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,524.70 C 1098.24,531.00 1098.24,539.40 1110.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,524.70 C 1098.24,531.00 1098.24,539.40 1110.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,524.70 C 1158.24,531.00 1158.24,539.40 1170.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,524.70 C 1158.24,531.00 1158.24,539.40 1170.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,524.70 C 1158.24,531.00 1158.24,539.40 1170.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,524.70 C 1218.24,531.00 1218.24,539.40 1230.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,524.70 C 1218.24,531.00 1218.24,539.40 1230.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,524.70 C 1218.24,531.00 1218.24,539.40 1230.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,524.70 C 1278.24,531.00 1278.24,539.40 1290.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,524.70 C 1278.24,531.00 1278.24,539.40 1290.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,524.70 C 1278.24,531.00 1278.24,539.40 1290.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,524.70 C 1338.24,531.00 1338.24,539.40 1350.00,545.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,524.70 C 1338.24,531.00 1338.24,539.40 1350.00,545.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,524.70 C 1338.24,531.00 1338.24,539.40 1350.00,545.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,584.70 C 138.24,591.00 138.24,599.40 150.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,584.70 C 138.24,591.00 138.24,599.40 150.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,584.70 C 138.24,591.00 138.24,599.40 150.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,584.70 C 198.24,591.00 198.24,599.40 210.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,584.70 C 198.24,591.00 198.24,599.40 210.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,584.70 C 198.24,591.00 198.24,599.40 210.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,584.70 C 258.24,591.00 258.24,599.40 270.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,584.70 C 258.24,591.00 258.24,599.40 270.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,584.70 C 258.24,591.00 258.24,599.40 270.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,584.70 C 318.24,591.00 318.24,599.40 330.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,584.70 C 318.24,591.00 318.24,599.40 330.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,584.70 C 318.24,591.00 318.24,599.40 330.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,584.70 C 378.24,591.00 378.24,599.40 390.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,584.70 C 378.24,591.00 378.24,599.40 390.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,584.70 C 378.24,591.00 378.24,599.40 390.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,584.70 C 438.24,591.00 438.24,599.40 450.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,584.70 C 438.24,591.00 438.24,599.40 450.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,584.70 C 438.24,591.00 438.24,599.40 450.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,584.70 C 498.24,591.00 498.24,599.40 510.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,584.70 C 498.24,591.00 498.24,599.40 510.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,584.70 C 498.24,591.00 498.24,599.40 510.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,584.70 C 558.24,591.00 558.24,599.40 570.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,584.70 C 558.24,591.00 558.24,599.40 570.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,584.70 C 558.24,591.00 558.24,599.40 570.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,584.70 C 618.24,591.00 618.24,599.40 630.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,584.70 C 618.24,591.00 618.24,599.40 630.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,584.70 C 618.24,591.00 618.24,599.40 630.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,584.70 C 678.24,591.00 678.24,599.40 690.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,584.70 C 678.24,591.00 678.24,599.40 690.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,584.70 C 678.24,591.00 678.24,599.40 690.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,584.70 C 738.24,591.00 738.24,599.40 750.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,584.70 C 738.24,591.00 738.24,599.40 750.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,584.70 C 738.24,591.00 738.24,599.40 750.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,584.70 C 798.24,591.00 798.24,599.40 810.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,584.70 C 798.24,591.00 798.24,599.40 810.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,584.70 C 798.24,591.00 798.24,599.40 810.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,584.70 C 858.24,591.00 858.24,599.40 870.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,584.70 C 858.24,591.00 858.24,599.40 870.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,584.70 C 858.24,591.00 858.24,599.40 870.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,584.70 C 918.24,591.00 918.24,599.40 930.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,584.70 C 918.24,591.00 918.24,599.40 930.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,584.70 C 918.24,591.00 918.24,599.40 930.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,584.70 C 978.24,591.00 978.24,599.40 990.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,584.70 C 978.24,591.00 978.24,599.40 990.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,584.70 C 978.24,591.00 978.24,599.40 990.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,584.70 C 1038.24,591.00 1038.24,599.40 1050.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,584.70 C 1038.24,591.00 1038.24,599.40 1050.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,584.70 C 1038.24,591.00 1038.24,599.40 1050.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,584.70 C 1098.24,591.00 1098.24,599.40 1110.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,584.70 C 1098.24,591.00 1098.24,599.40 1110.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,584.70 C 1098.24,591.00 1098.24,599.40 1110.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,584.70 C 1158.24,591.00 1158.24,599.40 1170.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,584.70 C 1158.24,591.00 1158.24,599.40 1170.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,584.70 C 1158.24,591.00 1158.24,599.40 1170.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,584.70 C 1218.24,591.00 1218.24,599.40 1230.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,584.70 C 1218.24,591.00 1218.24,599.40 1230.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,584.70 C 1218.24,591.00 1218.24,599.40 1230.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,584.70 C 1278.24,591.00 1278.24,599.40 1290.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,584.70 C 1278.24,591.00 1278.24,599.40 1290.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,584.70 C 1278.24,591.00 1278.24,599.40 1290.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,584.70 C 1338.24,591.00 1338.24,599.40 1350.00,605.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,584.70 C 1338.24,591.00 1338.24,599.40 1350.00,605.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,584.70 C 1338.24,591.00 1338.24,599.40 1350.00,605.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,644.70 C 138.24,651.00 138.24,659.40 150.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,644.70 C 138.24,651.00 138.24,659.40 150.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,644.70 C 138.24,651.00 138.24,659.40 150.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,644.70 C 198.24,651.00 198.24,659.40 210.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,644.70 C 198.24,651.00 198.24,659.40 210.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,644.70 C 198.24,651.00 198.24,659.40 210.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,644.70 C 258.24,651.00 258.24,659.40 270.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,644.70 C 258.24,651.00 258.24,659.40 270.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,644.70 C 258.24,651.00 258.24,659.40 270.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,644.70 C 318.24,651.00 318.24,659.40 330.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,644.70 C 318.24,651.00 318.24,659.40 330.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,644.70 C 318.24,651.00 318.24,659.40 330.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,644.70 C 378.24,651.00 378.24,659.40 390.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,644.70 C 378.24,651.00 378.24,659.40 390.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,644.70 C 378.24,651.00 378.24,659.40 390.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,644.70 C 438.24,651.00 438.24,659.40 450.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,644.70 C 438.24,651.00 438.24,659.40 450.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,644.70 C 438.24,651.00 438.24,659.40 450.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,644.70 C 498.24,651.00 498.24,659.40 510.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,644.70 C 498.24,651.00 498.24,659.40 510.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,644.70 C 498.24,651.00 498.24,659.40 510.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,644.70 C 558.24,651.00 558.24,659.40 570.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,644.70 C 558.24,651.00 558.24,659.40 570.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,644.70 C 558.24,651.00 558.24,659.40 570.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,644.70 C 618.24,651.00 618.24,659.40 630.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,644.70 C 618.24,651.00 618.24,659.40 630.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,644.70 C 618.24,651.00 618.24,659.40 630.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,644.70 C 678.24,651.00 678.24,659.40 690.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,644.70 C 678.24,651.00 678.24,659.40 690.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,644.70 C 678.24,651.00 678.24,659.40 690.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,644.70 C 738.24,651.00 738.24,659.40 750.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,644.70 C 738.24,651.00 738.24,659.40 750.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,644.70 C 738.24,651.00 738.24,659.40 750.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,644.70 C 798.24,651.00 798.24,659.40 810.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,644.70 C 798.24,651.00 798.24,659.40 810.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,644.70 C 798.24,651.00 798.24,659.40 810.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,644.70 C 858.24,651.00 858.24,659.40 870.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,644.70 C 858.24,651.00 858.24,659.40 870.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,644.70 C 858.24,651.00 858.24,659.40 870.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,644.70 C 918.24,651.00 918.24,659.40 930.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,644.70 C 918.24,651.00 918.24,659.40 930.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,644.70 C 918.24,651.00 918.24,659.40 930.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,644.70 C 978.24,651.00 978.24,659.40 990.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,644.70 C 978.24,651.00 978.24,659.40 990.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,644.70 C 978.24,651.00 978.24,659.40 990.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,644.70 C 1038.24,651.00 1038.24,659.40 1050.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,644.70 C 1038.24,651.00 1038.24,659.40 1050.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,644.70 C 1038.24,651.00 1038.24,659.40 1050.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,644.70 C 1098.24,651.00 1098.24,659.40 1110.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,644.70 C 1098.24,651.00 1098.24,659.40 1110.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,644.70 C 1098.24,651.00 1098.24,659.40 1110.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,644.70 C 1158.24,651.00 1158.24,659.40 1170.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,644.70 C 1158.24,651.00 1158.24,659.40 1170.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,644.70 C 1158.24,651.00 1158.24,659.40 1170.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,644.70 C 1218.24,651.00 1218.24,659.40 1230.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,644.70 C 1218.24,651.00 1218.24,659.40 1230.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,644.70 C 1218.24,651.00 1218.24,659.40 1230.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,644.70 C 1278.24,651.00 1278.24,659.40 1290.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,644.70 C 1278.24,651.00 1278.24,659.40 1290.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,644.70 C 1278.24,651.00 1278.24,659.40 1290.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,644.70 C 1338.24,651.00 1338.24,659.40 1350.00,665.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,644.70 C 1338.24,651.00 1338.24,659.40 1350.00,665.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,644.70 C 1338.24,651.00 1338.24,659.40 1350.00,665.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,704.70 C 138.24,711.00 138.24,719.40 150.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,704.70 C 138.24,711.00 138.24,719.40 150.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,704.70 C 138.24,711.00 138.24,719.40 150.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,704.70 C 198.24,711.00 198.24,719.40 210.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,704.70 C 198.24,711.00 198.24,719.40 210.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,704.70 C 198.24,711.00 198.24,719.40 210.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,704.70 C 258.24,711.00 258.24,719.40 270.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,704.70 C 258.24,711.00 258.24,719.40 270.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,704.70 C 258.24,711.00 258.24,719.40 270.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,704.70 C 318.24,711.00 318.24,719.40 330.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,704.70 C 318.24,711.00 318.24,719.40 330.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,704.70 C 318.24,711.00 318.24,719.40 330.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,704.70 C 378.24,711.00 378.24,719.40 390.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,704.70 C 378.24,711.00 378.24,719.40 390.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,704.70 C 378.24,711.00 378.24,719.40 390.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,704.70 C 438.24,711.00 438.24,719.40 450.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,704.70 C 438.24,711.00 438.24,719.40 450.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,704.70 C 438.24,711.00 438.24,719.40 450.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,704.70 C 498.24,711.00 498.24,719.40 510.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,704.70 C 498.24,711.00 498.24,719.40 510.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,704.70 C 498.24,711.00 498.24,719.40 510.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,704.70 C 558.24,711.00 558.24,719.40 570.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,704.70 C 558.24,711.00 558.24,719.40 570.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,704.70 C 558.24,711.00 558.24,719.40 570.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,704.70 C 618.24,711.00 618.24,719.40 630.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,704.70 C 618.24,711.00 618.24,719.40 630.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,704.70 C 618.24,711.00 618.24,719.40 630.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,704.70 C 678.24,711.00 678.24,719.40 690.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,704.70 C 678.24,711.00 678.24,719.40 690.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,704.70 C 678.24,711.00 678.24,719.40 690.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,704.70 C 738.24,711.00 738.24,719.40 750.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,704.70 C 738.24,711.00 738.24,719.40 750.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,704.70 C 738.24,711.00 738.24,719.40 750.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,704.70 C 798.24,711.00 798.24,719.40 810.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,704.70 C 798.24,711.00 798.24,719.40 810.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,704.70 C 798.24,711.00 798.24,719.40 810.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,704.70 C 858.24,711.00 858.24,719.40 870.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,704.70 C 858.24,711.00 858.24,719.40 870.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,704.70 C 858.24,711.00 858.24,719.40 870.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,704.70 C 918.24,711.00 918.24,719.40 930.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,704.70 C 918.24,711.00 918.24,719.40 930.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,704.70 C 918.24,711.00 918.24,719.40 930.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,704.70 C 978.24,711.00 978.24,719.40 990.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,704.70 C 978.24,711.00 978.24,719.40 990.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,704.70 C 978.24,711.00 978.24,719.40 990.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,704.70 C 1038.24,711.00 1038.24,719.40 1050.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,704.70 C 1038.24,711.00 1038.24,719.40 1050.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,704.70 C 1038.24,711.00 1038.24,719.40 1050.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,704.70 C 1098.24,711.00 1098.24,719.40 1110.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,704.70 C 1098.24,711.00 1098.24,719.40 1110.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,704.70 C 1098.24,711.00 1098.24,719.40 1110.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,704.70 C 1158.24,711.00 1158.24,719.40 1170.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,704.70 C 1158.24,711.00 1158.24,719.40 1170.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,704.70 C 1158.24,711.00 1158.24,719.40 1170.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,704.70 C 1218.24,711.00 1218.24,719.40 1230.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,704.70 C 1218.24,711.00 1218.24,719.40 1230.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,704.70 C 1218.24,711.00 1218.24,719.40 1230.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,704.70 C 1278.24,711.00 1278.24,719.40 1290.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,704.70 C 1278.24,711.00 1278.24,719.40 1290.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,704.70 C 1278.24,711.00 1278.24,719.40 1290.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,704.70 C 1338.24,711.00 1338.24,719.40 1350.00,725.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,704.70 C 1338.24,711.00 1338.24,719.40 1350.00,725.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,704.70 C 1338.24,711.00 1338.24,719.40 1350.00,725.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,764.70 C 138.24,771.00 138.24,779.40 150.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,764.70 C 138.24,771.00 138.24,779.40 150.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,764.70 C 138.24,771.00 138.24,779.40 150.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,764.70 C 198.24,771.00 198.24,779.40 210.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,764.70 C 198.24,771.00 198.24,779.40 210.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,764.70 C 198.24,771.00 198.24,779.40 210.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,764.70 C 258.24,771.00 258.24,779.40 270.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,764.70 C 258.24,771.00 258.24,779.40 270.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,764.70 C 258.24,771.00 258.24,779.40 270.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,764.70 C 318.24,771.00 318.24,779.40 330.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,764.70 C 318.24,771.00 318.24,779.40 330.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,764.70 C 318.24,771.00 318.24,779.40 330.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,764.70 C 378.24,771.00 378.24,779.40 390.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,764.70 C 378.24,771.00 378.24,779.40 390.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,764.70 C 378.24,771.00 378.24,779.40 390.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,764.70 C 438.24,771.00 438.24,779.40 450.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,764.70 C 438.24,771.00 438.24,779.40 450.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,764.70 C 438.24,771.00 438.24,779.40 450.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,764.70 C 498.24,771.00 498.24,779.40 510.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,764.70 C 498.24,771.00 498.24,779.40 510.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,764.70 C 498.24,771.00 498.24,779.40 510.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,764.70 C 558.24,771.00 558.24,779.40 570.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,764.70 C 558.24,771.00 558.24,779.40 570.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,764.70 C 558.24,771.00 558.24,779.40 570.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,764.70 C 618.24,771.00 618.24,779.40 630.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,764.70 C 618.24,771.00 618.24,779.40 630.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,764.70 C 618.24,771.00 618.24,779.40 630.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,764.70 C 678.24,771.00 678.24,779.40 690.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,764.70 C 678.24,771.00 678.24,779.40 690.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,764.70 C 678.24,771.00 678.24,779.40 690.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,764.70 C 738.24,771.00 738.24,779.40 750.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,764.70 C 738.24,771.00 738.24,779.40 750.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,764.70 C 738.24,771.00 738.24,779.40 750.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,764.70 C 798.24,771.00 798.24,779.40 810.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,764.70 C 798.24,771.00 798.24,779.40 810.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,764.70 C 798.24,771.00 798.24,779.40 810.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,764.70 C 858.24,771.00 858.24,779.40 870.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,764.70 C 858.24,771.00 858.24,779.40 870.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,764.70 C 858.24,771.00 858.24,779.40 870.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,764.70 C 918.24,771.00 918.24,779.40 930.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,764.70 C 918.24,771.00 918.24,779.40 930.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,764.70 C 918.24,771.00 918.24,779.40 930.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,764.70 C 978.24,771.00 978.24,779.40 990.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,764.70 C 978.24,771.00 978.24,779.40 990.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,764.70 C 978.24,771.00 978.24,779.40 990.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,764.70 C 1038.24,771.00 1038.24,779.40 1050.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,764.70 C 1038.24,771.00 1038.24,779.40 1050.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,764.70 C 1038.24,771.00 1038.24,779.40 1050.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,764.70 C 1098.24,771.00 1098.24,779.40 1110.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,764.70 C 1098.24,771.00 1098.24,779.40 1110.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,764.70 C 1098.24,771.00 1098.24,779.40 1110.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,764.70 C 1158.24,771.00 1158.24,779.40 1170.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,764.70 C 1158.24,771.00 1158.24,779.40 1170.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,764.70 C 1158.24,771.00 1158.24,779.40 1170.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,764.70 C 1218.24,771.00 1218.24,779.40 1230.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,764.70 C 1218.24,771.00 1218.24,779.40 1230.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,764.70 C 1218.24,771.00 1218.24,779.40 1230.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,764.70 C 1278.24,771.00 1278.24,779.40 1290.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,764.70 C 1278.24,771.00 1278.24,779.40 1290.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,764.70 C 1278.24,771.00 1278.24,779.40 1290.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,764.70 C 1338.24,771.00 1338.24,779.40 1350.00,785.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,764.70 C 1338.24,771.00 1338.24,779.40 1350.00,785.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,764.70 C 1338.24,771.00 1338.24,779.40 1350.00,785.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,824.70 C 138.24,831.00 138.24,839.40 150.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,824.70 C 138.24,831.00 138.24,839.40 150.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,824.70 C 138.24,831.00 138.24,839.40 150.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,824.70 C 198.24,831.00 198.24,839.40 210.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,824.70 C 198.24,831.00 198.24,839.40 210.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,824.70 C 198.24,831.00 198.24,839.40 210.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,824.70 C 258.24,831.00 258.24,839.40 270.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,824.70 C 258.24,831.00 258.24,839.40 270.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,824.70 C 258.24,831.00 258.24,839.40 270.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,824.70 C 318.24,831.00 318.24,839.40 330.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,824.70 C 318.24,831.00 318.24,839.40 330.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,824.70 C 318.24,831.00 318.24,839.40 330.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,824.70 C 378.24,831.00 378.24,839.40 390.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,824.70 C 378.24,831.00 378.24,839.40 390.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,824.70 C 378.24,831.00 378.24,839.40 390.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,824.70 C 438.24,831.00 438.24,839.40 450.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,824.70 C 438.24,831.00 438.24,839.40 450.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,824.70 C 438.24,831.00 438.24,839.40 450.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,824.70 C 498.24,831.00 498.24,839.40 510.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,824.70 C 498.24,831.00 498.24,839.40 510.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,824.70 C 498.24,831.00 498.24,839.40 510.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,824.70 C 558.24,831.00 558.24,839.40 570.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,824.70 C 558.24,831.00 558.24,839.40 570.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,824.70 C 558.24,831.00 558.24,839.40 570.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,824.70 C 618.24,831.00 618.24,839.40 630.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,824.70 C 618.24,831.00 618.24,839.40 630.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,824.70 C 618.24,831.00 618.24,839.40 630.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,824.70 C 678.24,831.00 678.24,839.40 690.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,824.70 C 678.24,831.00 678.24,839.40 690.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,824.70 C 678.24,831.00 678.24,839.40 690.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,824.70 C 738.24,831.00 738.24,839.40 750.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,824.70 C 738.24,831.00 738.24,839.40 750.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,824.70 C 738.24,831.00 738.24,839.40 750.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,824.70 C 798.24,831.00 798.24,839.40 810.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,824.70 C 798.24,831.00 798.24,839.40 810.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,824.70 C 798.24,831.00 798.24,839.40 810.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,824.70 C 858.24,831.00 858.24,839.40 870.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,824.70 C 858.24,831.00 858.24,839.40 870.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,824.70 C 858.24,831.00 858.24,839.40 870.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,824.70 C 918.24,831.00 918.24,839.40 930.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,824.70 C 918.24,831.00 918.24,839.40 930.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,824.70 C 918.24,831.00 918.24,839.40 930.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,824.70 C 978.24,831.00 978.24,839.40 990.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,824.70 C 978.24,831.00 978.24,839.40 990.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,824.70 C 978.24,831.00 978.24,839.40 990.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,824.70 C 1038.24,831.00 1038.24,839.40 1050.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,824.70 C 1038.24,831.00 1038.24,839.40 1050.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,824.70 C 1038.24,831.00 1038.24,839.40 1050.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,824.70 C 1098.24,831.00 1098.24,839.40 1110.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,824.70 C 1098.24,831.00 1098.24,839.40 1110.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,824.70 C 1098.24,831.00 1098.24,839.40 1110.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,824.70 C 1158.24,831.00 1158.24,839.40 1170.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,824.70 C 1158.24,831.00 1158.24,839.40 1170.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,824.70 C 1158.24,831.00 1158.24,839.40 1170.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,824.70 C 1218.24,831.00 1218.24,839.40 1230.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,824.70 C 1218.24,831.00 1218.24,839.40 1230.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,824.70 C 1218.24,831.00 1218.24,839.40 1230.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,824.70 C 1278.24,831.00 1278.24,839.40 1290.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,824.70 C 1278.24,831.00 1278.24,839.40 1290.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,824.70 C 1278.24,831.00 1278.24,839.40 1290.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,824.70 C 1338.24,831.00 1338.24,839.40 1350.00,845.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,824.70 C 1338.24,831.00 1338.24,839.40 1350.00,845.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,824.70 C 1338.24,831.00 1338.24,839.40 1350.00,845.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,884.70 C 138.24,891.00 138.24,899.40 150.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,884.70 C 138.24,891.00 138.24,899.40 150.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,884.70 C 138.24,891.00 138.24,899.40 150.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,884.70 C 198.24,891.00 198.24,899.40 210.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,884.70 C 198.24,891.00 198.24,899.40 210.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,884.70 C 198.24,891.00 198.24,899.40 210.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,884.70 C 258.24,891.00 258.24,899.40 270.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,884.70 C 258.24,891.00 258.24,899.40 270.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,884.70 C 258.24,891.00 258.24,899.40 270.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,884.70 C 318.24,891.00 318.24,899.40 330.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,884.70 C 318.24,891.00 318.24,899.40 330.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,884.70 C 318.24,891.00 318.24,899.40 330.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,884.70 C 378.24,891.00 378.24,899.40 390.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,884.70 C 378.24,891.00 378.24,899.40 390.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,884.70 C 378.24,891.00 378.24,899.40 390.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,884.70 C 438.24,891.00 438.24,899.40 450.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,884.70 C 438.24,891.00 438.24,899.40 450.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,884.70 C 438.24,891.00 438.24,899.40 450.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,884.70 C 498.24,891.00 498.24,899.40 510.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,884.70 C 498.24,891.00 498.24,899.40 510.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,884.70 C 498.24,891.00 498.24,899.40 510.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,884.70 C 558.24,891.00 558.24,899.40 570.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,884.70 C 558.24,891.00 558.24,899.40 570.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,884.70 C 558.24,891.00 558.24,899.40 570.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,884.70 C 618.24,891.00 618.24,899.40 630.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,884.70 C 618.24,891.00 618.24,899.40 630.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,884.70 C 618.24,891.00 618.24,899.40 630.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,884.70 C 678.24,891.00 678.24,899.40 690.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,884.70 C 678.24,891.00 678.24,899.40 690.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,884.70 C 678.24,891.00 678.24,899.40 690.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,884.70 C 738.24,891.00 738.24,899.40 750.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,884.70 C 738.24,891.00 738.24,899.40 750.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,884.70 C 738.24,891.00 738.24,899.40 750.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,884.70 C 798.24,891.00 798.24,899.40 810.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,884.70 C 798.24,891.00 798.24,899.40 810.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,884.70 C 798.24,891.00 798.24,899.40 810.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,884.70 C 858.24,891.00 858.24,899.40 870.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,884.70 C 858.24,891.00 858.24,899.40 870.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,884.70 C 858.24,891.00 858.24,899.40 870.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,884.70 C 918.24,891.00 918.24,899.40 930.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,884.70 C 918.24,891.00 918.24,899.40 930.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,884.70 C 918.24,891.00 918.24,899.40 930.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,884.70 C 978.24,891.00 978.24,899.40 990.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,884.70 C 978.24,891.00 978.24,899.40 990.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,884.70 C 978.24,891.00 978.24,899.40 990.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,884.70 C 1038.24,891.00 1038.24,899.40 1050.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,884.70 C 1038.24,891.00 1038.24,899.40 1050.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,884.70 C 1038.24,891.00 1038.24,899.40 1050.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,884.70 C 1098.24,891.00 1098.24,899.40 1110.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,884.70 C 1098.24,891.00 1098.24,899.40 1110.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,884.70 C 1098.24,891.00 1098.24,899.40 1110.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,884.70 C 1158.24,891.00 1158.24,899.40 1170.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,884.70 C 1158.24,891.00 1158.24,899.40 1170.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,884.70 C 1158.24,891.00 1158.24,899.40 1170.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,884.70 C 1218.24,891.00 1218.24,899.40 1230.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,884.70 C 1218.24,891.00 1218.24,899.40 1230.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,884.70 C 1218.24,891.00 1218.24,899.40 1230.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,884.70 C 1278.24,891.00 1278.24,899.40 1290.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,884.70 C 1278.24,891.00 1278.24,899.40 1290.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,884.70 C 1278.24,891.00 1278.24,899.40 1290.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,884.70 C 1338.24,891.00 1338.24,899.40 1350.00,905.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,884.70 C 1338.24,891.00 1338.24,899.40 1350.00,905.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,884.70 C 1338.24,891.00 1338.24,899.40 1350.00,905.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,944.70 C 138.24,951.00 138.24,959.40 150.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,944.70 C 138.24,951.00 138.24,959.40 150.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,944.70 C 138.24,951.00 138.24,959.40 150.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,944.70 C 198.24,951.00 198.24,959.40 210.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,944.70 C 198.24,951.00 198.24,959.40 210.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,944.70 C 198.24,951.00 198.24,959.40 210.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,944.70 C 258.24,951.00 258.24,959.40 270.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,944.70 C 258.24,951.00 258.24,959.40 270.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,944.70 C 258.24,951.00 258.24,959.40 270.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,944.70 C 318.24,951.00 318.24,959.40 330.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,944.70 C 318.24,951.00 318.24,959.40 330.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,944.70 C 318.24,951.00 318.24,959.40 330.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,944.70 C 378.24,951.00 378.24,959.40 390.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,944.70 C 378.24,951.00 378.24,959.40 390.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,944.70 C 378.24,951.00 378.24,959.40 390.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,944.70 C 438.24,951.00 438.24,959.40 450.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,944.70 C 438.24,951.00 438.24,959.40 450.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,944.70 C 438.24,951.00 438.24,959.40 450.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,944.70 C 498.24,951.00 498.24,959.40 510.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,944.70 C 498.24,951.00 498.24,959.40 510.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,944.70 C 498.24,951.00 498.24,959.40 510.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,944.70 C 558.24,951.00 558.24,959.40 570.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,944.70 C 558.24,951.00 558.24,959.40 570.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,944.70 C 558.24,951.00 558.24,959.40 570.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,944.70 C 618.24,951.00 618.24,959.40 630.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,944.70 C 618.24,951.00 618.24,959.40 630.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,944.70 C 618.24,951.00 618.24,959.40 630.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,944.70 C 678.24,951.00 678.24,959.40 690.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,944.70 C 678.24,951.00 678.24,959.40 690.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,944.70 C 678.24,951.00 678.24,959.40 690.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,944.70 C 738.24,951.00 738.24,959.40 750.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,944.70 C 738.24,951.00 738.24,959.40 750.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,944.70 C 738.24,951.00 738.24,959.40 750.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,944.70 C 798.24,951.00 798.24,959.40 810.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,944.70 C 798.24,951.00 798.24,959.40 810.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,944.70 C 798.24,951.00 798.24,959.40 810.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,944.70 C 858.24,951.00 858.24,959.40 870.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,944.70 C 858.24,951.00 858.24,959.40 870.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,944.70 C 858.24,951.00 858.24,959.40 870.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,944.70 C 918.24,951.00 918.24,959.40 930.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,944.70 C 918.24,951.00 918.24,959.40 930.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,944.70 C 918.24,951.00 918.24,959.40 930.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,944.70 C 978.24,951.00 978.24,959.40 990.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,944.70 C 978.24,951.00 978.24,959.40 990.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,944.70 C 978.24,951.00 978.24,959.40 990.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,944.70 C 1038.24,951.00 1038.24,959.40 1050.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,944.70 C 1038.24,951.00 1038.24,959.40 1050.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,944.70 C 1038.24,951.00 1038.24,959.40 1050.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,944.70 C 1098.24,951.00 1098.24,959.40 1110.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,944.70 C 1098.24,951.00 1098.24,959.40 1110.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,944.70 C 1098.24,951.00 1098.24,959.40 1110.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,944.70 C 1158.24,951.00 1158.24,959.40 1170.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,944.70 C 1158.24,951.00 1158.24,959.40 1170.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,944.70 C 1158.24,951.00 1158.24,959.40 1170.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,944.70 C 1218.24,951.00 1218.24,959.40 1230.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,944.70 C 1218.24,951.00 1218.24,959.40 1230.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,944.70 C 1218.24,951.00 1218.24,959.40 1230.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,944.70 C 1278.24,951.00 1278.24,959.40 1290.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,944.70 C 1278.24,951.00 1278.24,959.40 1290.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,944.70 C 1278.24,951.00 1278.24,959.40 1290.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,944.70 C 1338.24,951.00 1338.24,959.40 1350.00,965.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,944.70 C 1338.24,951.00 1338.24,959.40 1350.00,965.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,944.70 C 1338.24,951.00 1338.24,959.40 1350.00,965.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,1004.70 C 138.24,1011.00 138.24,1019.40 150.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,1004.70 C 138.24,1011.00 138.24,1019.40 150.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,1004.70 C 138.24,1011.00 138.24,1019.40 150.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,1004.70 C 198.24,1011.00 198.24,1019.40 210.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,1004.70 C 198.24,1011.00 198.24,1019.40 210.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,1004.70 C 198.24,1011.00 198.24,1019.40 210.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,1004.70 C 258.24,1011.00 258.24,1019.40 270.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,1004.70 C 258.24,1011.00 258.24,1019.40 270.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,1004.70 C 258.24,1011.00 258.24,1019.40 270.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,1004.70 C 318.24,1011.00 318.24,1019.40 330.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,1004.70 C 318.24,1011.00 318.24,1019.40 330.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,1004.70 C 318.24,1011.00 318.24,1019.40 330.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,1004.70 C 378.24,1011.00 378.24,1019.40 390.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,1004.70 C 378.24,1011.00 378.24,1019.40 390.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,1004.70 C 378.24,1011.00 378.24,1019.40 390.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,1004.70 C 438.24,1011.00 438.24,1019.40 450.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,1004.70 C 438.24,1011.00 438.24,1019.40 450.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,1004.70 C 438.24,1011.00 438.24,1019.40 450.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,1004.70 C 498.24,1011.00 498.24,1019.40 510.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,1004.70 C 498.24,1011.00 498.24,1019.40 510.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,1004.70 C 498.24,1011.00 498.24,1019.40 510.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,1004.70 C 558.24,1011.00 558.24,1019.40 570.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,1004.70 C 558.24,1011.00 558.24,1019.40 570.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,1004.70 C 558.24,1011.00 558.24,1019.40 570.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,1004.70 C 618.24,1011.00 618.24,1019.40 630.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,1004.70 C 618.24,1011.00 618.24,1019.40 630.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,1004.70 C 618.24,1011.00 618.24,1019.40 630.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,1004.70 C 678.24,1011.00 678.24,1019.40 690.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,1004.70 C 678.24,1011.00 678.24,1019.40 690.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,1004.70 C 678.24,1011.00 678.24,1019.40 690.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,1004.70 C 738.24,1011.00 738.24,1019.40 750.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,1004.70 C 738.24,1011.00 738.24,1019.40 750.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,1004.70 C 738.24,1011.00 738.24,1019.40 750.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,1004.70 C 798.24,1011.00 798.24,1019.40 810.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,1004.70 C 798.24,1011.00 798.24,1019.40 810.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,1004.70 C 798.24,1011.00 798.24,1019.40 810.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,1004.70 C 858.24,1011.00 858.24,1019.40 870.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,1004.70 C 858.24,1011.00 858.24,1019.40 870.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,1004.70 C 858.24,1011.00 858.24,1019.40 870.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,1004.70 C 918.24,1011.00 918.24,1019.40 930.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,1004.70 C 918.24,1011.00 918.24,1019.40 930.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,1004.70 C 918.24,1011.00 918.24,1019.40 930.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,1004.70 C 978.24,1011.00 978.24,1019.40 990.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,1004.70 C 978.24,1011.00 978.24,1019.40 990.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,1004.70 C 978.24,1011.00 978.24,1019.40 990.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,1004.70 C 1038.24,1011.00 1038.24,1019.40 1050.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,1004.70 C 1038.24,1011.00 1038.24,1019.40 1050.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,1004.70 C 1038.24,1011.00 1038.24,1019.40 1050.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,1004.70 C 1098.24,1011.00 1098.24,1019.40 1110.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,1004.70 C 1098.24,1011.00 1098.24,1019.40 1110.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,1004.70 C 1098.24,1011.00 1098.24,1019.40 1110.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,1004.70 C 1158.24,1011.00 1158.24,1019.40 1170.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,1004.70 C 1158.24,1011.00 1158.24,1019.40 1170.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,1004.70 C 1158.24,1011.00 1158.24,1019.40 1170.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,1004.70 C 1218.24,1011.00 1218.24,1019.40 1230.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,1004.70 C 1218.24,1011.00 1218.24,1019.40 1230.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,1004.70 C 1218.24,1011.00 1218.24,1019.40 1230.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,1004.70 C 1278.24,1011.00 1278.24,1019.40 1290.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,1004.70 C 1278.24,1011.00 1278.24,1019.40 1290.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,1004.70 C 1278.24,1011.00 1278.24,1019.40 1290.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,1004.70 C 1338.24,1011.00 1338.24,1019.40 1350.00,1025.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,1004.70 C 1338.24,1011.00 1338.24,1019.40 1350.00,1025.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,1004.70 C 1338.24,1011.00 1338.24,1019.40 1350.00,1025.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,1064.70 C 138.24,1071.00 138.24,1079.40 150.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,1064.70 C 138.24,1071.00 138.24,1079.40 150.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,1064.70 C 138.24,1071.00 138.24,1079.40 150.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,1064.70 C 198.24,1071.00 198.24,1079.40 210.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,1064.70 C 198.24,1071.00 198.24,1079.40 210.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,1064.70 C 198.24,1071.00 198.24,1079.40 210.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,1064.70 C 258.24,1071.00 258.24,1079.40 270.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,1064.70 C 258.24,1071.00 258.24,1079.40 270.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,1064.70 C 258.24,1071.00 258.24,1079.40 270.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,1064.70 C 318.24,1071.00 318.24,1079.40 330.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,1064.70 C 318.24,1071.00 318.24,1079.40 330.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,1064.70 C 318.24,1071.00 318.24,1079.40 330.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,1064.70 C 378.24,1071.00 378.24,1079.40 390.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,1064.70 C 378.24,1071.00 378.24,1079.40 390.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,1064.70 C 378.24,1071.00 378.24,1079.40 390.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,1064.70 C 438.24,1071.00 438.24,1079.40 450.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,1064.70 C 438.24,1071.00 438.24,1079.40 450.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,1064.70 C 438.24,1071.00 438.24,1079.40 450.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,1064.70 C 498.24,1071.00 498.24,1079.40 510.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,1064.70 C 498.24,1071.00 498.24,1079.40 510.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,1064.70 C 498.24,1071.00 498.24,1079.40 510.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,1064.70 C 558.24,1071.00 558.24,1079.40 570.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,1064.70 C 558.24,1071.00 558.24,1079.40 570.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,1064.70 C 558.24,1071.00 558.24,1079.40 570.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,1064.70 C 618.24,1071.00 618.24,1079.40 630.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,1064.70 C 618.24,1071.00 618.24,1079.40 630.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,1064.70 C 618.24,1071.00 618.24,1079.40 630.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,1064.70 C 678.24,1071.00 678.24,1079.40 690.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,1064.70 C 678.24,1071.00 678.24,1079.40 690.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,1064.70 C 678.24,1071.00 678.24,1079.40 690.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,1064.70 C 738.24,1071.00 738.24,1079.40 750.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,1064.70 C 738.24,1071.00 738.24,1079.40 750.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,1064.70 C 738.24,1071.00 738.24,1079.40 750.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,1064.70 C 798.24,1071.00 798.24,1079.40 810.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,1064.70 C 798.24,1071.00 798.24,1079.40 810.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,1064.70 C 798.24,1071.00 798.24,1079.40 810.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,1064.70 C 858.24,1071.00 858.24,1079.40 870.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,1064.70 C 858.24,1071.00 858.24,1079.40 870.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,1064.70 C 858.24,1071.00 858.24,1079.40 870.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,1064.70 C 918.24,1071.00 918.24,1079.40 930.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,1064.70 C 918.24,1071.00 918.24,1079.40 930.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,1064.70 C 918.24,1071.00 918.24,1079.40 930.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,1064.70 C 978.24,1071.00 978.24,1079.40 990.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,1064.70 C 978.24,1071.00 978.24,1079.40 990.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,1064.70 C 978.24,1071.00 978.24,1079.40 990.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,1064.70 C 1038.24,1071.00 1038.24,1079.40 1050.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,1064.70 C 1038.24,1071.00 1038.24,1079.40 1050.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,1064.70 C 1038.24,1071.00 1038.24,1079.40 1050.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,1064.70 C 1098.24,1071.00 1098.24,1079.40 1110.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,1064.70 C 1098.24,1071.00 1098.24,1079.40 1110.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,1064.70 C 1098.24,1071.00 1098.24,1079.40 1110.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,1064.70 C 1158.24,1071.00 1158.24,1079.40 1170.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,1064.70 C 1158.24,1071.00 1158.24,1079.40 1170.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,1064.70 C 1158.24,1071.00 1158.24,1079.40 1170.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,1064.70 C 1218.24,1071.00 1218.24,1079.40 1230.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,1064.70 C 1218.24,1071.00 1218.24,1079.40 1230.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,1064.70 C 1218.24,1071.00 1218.24,1079.40 1230.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,1064.70 C 1278.24,1071.00 1278.24,1079.40 1290.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,1064.70 C 1278.24,1071.00 1278.24,1079.40 1290.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,1064.70 C 1278.24,1071.00 1278.24,1079.40 1290.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,1064.70 C 1338.24,1071.00 1338.24,1079.40 1350.00,1085.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,1064.70 C 1338.24,1071.00 1338.24,1079.40 1350.00,1085.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,1064.70 C 1338.24,1071.00 1338.24,1079.40 1350.00,1085.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,1124.70 C 138.24,1131.00 138.24,1139.40 150.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,1124.70 C 138.24,1131.00 138.24,1139.40 150.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,1124.70 C 138.24,1131.00 138.24,1139.40 150.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,1124.70 C 198.24,1131.00 198.24,1139.40 210.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,1124.70 C 198.24,1131.00 198.24,1139.40 210.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,1124.70 C 198.24,1131.00 198.24,1139.40 210.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,1124.70 C 258.24,1131.00 258.24,1139.40 270.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,1124.70 C 258.24,1131.00 258.24,1139.40 270.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,1124.70 C 258.24,1131.00 258.24,1139.40 270.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,1124.70 C 318.24,1131.00 318.24,1139.40 330.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,1124.70 C 318.24,1131.00 318.24,1139.40 330.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,1124.70 C 318.24,1131.00 318.24,1139.40 330.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,1124.70 C 378.24,1131.00 378.24,1139.40 390.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,1124.70 C 378.24,1131.00 378.24,1139.40 390.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,1124.70 C 378.24,1131.00 378.24,1139.40 390.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,1124.70 C 438.24,1131.00 438.24,1139.40 450.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,1124.70 C 438.24,1131.00 438.24,1139.40 450.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,1124.70 C 438.24,1131.00 438.24,1139.40 450.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,1124.70 C 498.24,1131.00 498.24,1139.40 510.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,1124.70 C 498.24,1131.00 498.24,1139.40 510.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,1124.70 C 498.24,1131.00 498.24,1139.40 510.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,1124.70 C 558.24,1131.00 558.24,1139.40 570.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,1124.70 C 558.24,1131.00 558.24,1139.40 570.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,1124.70 C 558.24,1131.00 558.24,1139.40 570.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,1124.70 C 618.24,1131.00 618.24,1139.40 630.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,1124.70 C 618.24,1131.00 618.24,1139.40 630.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,1124.70 C 618.24,1131.00 618.24,1139.40 630.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,1124.70 C 678.24,1131.00 678.24,1139.40 690.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,1124.70 C 678.24,1131.00 678.24,1139.40 690.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,1124.70 C 678.24,1131.00 678.24,1139.40 690.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,1124.70 C 738.24,1131.00 738.24,1139.40 750.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,1124.70 C 738.24,1131.00 738.24,1139.40 750.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,1124.70 C 738.24,1131.00 738.24,1139.40 750.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,1124.70 C 798.24,1131.00 798.24,1139.40 810.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,1124.70 C 798.24,1131.00 798.24,1139.40 810.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,1124.70 C 798.24,1131.00 798.24,1139.40 810.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,1124.70 C 858.24,1131.00 858.24,1139.40 870.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,1124.70 C 858.24,1131.00 858.24,1139.40 870.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,1124.70 C 858.24,1131.00 858.24,1139.40 870.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,1124.70 C 918.24,1131.00 918.24,1139.40 930.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,1124.70 C 918.24,1131.00 918.24,1139.40 930.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,1124.70 C 918.24,1131.00 918.24,1139.40 930.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,1124.70 C 978.24,1131.00 978.24,1139.40 990.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,1124.70 C 978.24,1131.00 978.24,1139.40 990.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,1124.70 C 978.24,1131.00 978.24,1139.40 990.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,1124.70 C 1038.24,1131.00 1038.24,1139.40 1050.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,1124.70 C 1038.24,1131.00 1038.24,1139.40 1050.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,1124.70 C 1038.24,1131.00 1038.24,1139.40 1050.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,1124.70 C 1098.24,1131.00 1098.24,1139.40 1110.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,1124.70 C 1098.24,1131.00 1098.24,1139.40 1110.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,1124.70 C 1098.24,1131.00 1098.24,1139.40 1110.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,1124.70 C 1158.24,1131.00 1158.24,1139.40 1170.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,1124.70 C 1158.24,1131.00 1158.24,1139.40 1170.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,1124.70 C 1158.24,1131.00 1158.24,1139.40 1170.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,1124.70 C 1218.24,1131.00 1218.24,1139.40 1230.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,1124.70 C 1218.24,1131.00 1218.24,1139.40 1230.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,1124.70 C 1218.24,1131.00 1218.24,1139.40 1230.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,1124.70 C 1278.24,1131.00 1278.24,1139.40 1290.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,1124.70 C 1278.24,1131.00 1278.24,1139.40 1290.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,1124.70 C 1278.24,1131.00 1278.24,1139.40 1290.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,1124.70 C 1338.24,1131.00 1338.24,1139.40 1350.00,1145.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,1124.70 C 1338.24,1131.00 1338.24,1139.40 1350.00,1145.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,1124.70 C 1338.24,1131.00 1338.24,1139.40 1350.00,1145.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,1184.70 C 138.24,1191.00 138.24,1199.40 150.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,1184.70 C 138.24,1191.00 138.24,1199.40 150.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,1184.70 C 138.24,1191.00 138.24,1199.40 150.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,1184.70 C 198.24,1191.00 198.24,1199.40 210.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,1184.70 C 198.24,1191.00 198.24,1199.40 210.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,1184.70 C 198.24,1191.00 198.24,1199.40 210.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,1184.70 C 258.24,1191.00 258.24,1199.40 270.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,1184.70 C 258.24,1191.00 258.24,1199.40 270.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,1184.70 C 258.24,1191.00 258.24,1199.40 270.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,1184.70 C 318.24,1191.00 318.24,1199.40 330.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,1184.70 C 318.24,1191.00 318.24,1199.40 330.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,1184.70 C 318.24,1191.00 318.24,1199.40 330.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,1184.70 C 378.24,1191.00 378.24,1199.40 390.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,1184.70 C 378.24,1191.00 378.24,1199.40 390.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,1184.70 C 378.24,1191.00 378.24,1199.40 390.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,1184.70 C 438.24,1191.00 438.24,1199.40 450.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,1184.70 C 438.24,1191.00 438.24,1199.40 450.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,1184.70 C 438.24,1191.00 438.24,1199.40 450.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,1184.70 C 498.24,1191.00 498.24,1199.40 510.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,1184.70 C 498.24,1191.00 498.24,1199.40 510.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,1184.70 C 498.24,1191.00 498.24,1199.40 510.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,1184.70 C 558.24,1191.00 558.24,1199.40 570.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,1184.70 C 558.24,1191.00 558.24,1199.40 570.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,1184.70 C 558.24,1191.00 558.24,1199.40 570.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,1184.70 C 618.24,1191.00 618.24,1199.40 630.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,1184.70 C 618.24,1191.00 618.24,1199.40 630.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,1184.70 C 618.24,1191.00 618.24,1199.40 630.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,1184.70 C 678.24,1191.00 678.24,1199.40 690.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,1184.70 C 678.24,1191.00 678.24,1199.40 690.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,1184.70 C 678.24,1191.00 678.24,1199.40 690.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,1184.70 C 738.24,1191.00 738.24,1199.40 750.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,1184.70 C 738.24,1191.00 738.24,1199.40 750.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,1184.70 C 738.24,1191.00 738.24,1199.40 750.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,1184.70 C 798.24,1191.00 798.24,1199.40 810.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,1184.70 C 798.24,1191.00 798.24,1199.40 810.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,1184.70 C 798.24,1191.00 798.24,1199.40 810.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,1184.70 C 858.24,1191.00 858.24,1199.40 870.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,1184.70 C 858.24,1191.00 858.24,1199.40 870.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,1184.70 C 858.24,1191.00 858.24,1199.40 870.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,1184.70 C 918.24,1191.00 918.24,1199.40 930.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,1184.70 C 918.24,1191.00 918.24,1199.40 930.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,1184.70 C 918.24,1191.00 918.24,1199.40 930.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,1184.70 C 978.24,1191.00 978.24,1199.40 990.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,1184.70 C 978.24,1191.00 978.24,1199.40 990.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,1184.70 C 978.24,1191.00 978.24,1199.40 990.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,1184.70 C 1038.24,1191.00 1038.24,1199.40 1050.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,1184.70 C 1038.24,1191.00 1038.24,1199.40 1050.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,1184.70 C 1038.24,1191.00 1038.24,1199.40 1050.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,1184.70 C 1098.24,1191.00 1098.24,1199.40 1110.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,1184.70 C 1098.24,1191.00 1098.24,1199.40 1110.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,1184.70 C 1098.24,1191.00 1098.24,1199.40 1110.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,1184.70 C 1158.24,1191.00 1158.24,1199.40 1170.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,1184.70 C 1158.24,1191.00 1158.24,1199.40 1170.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,1184.70 C 1158.24,1191.00 1158.24,1199.40 1170.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,1184.70 C 1218.24,1191.00 1218.24,1199.40 1230.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,1184.70 C 1218.24,1191.00 1218.24,1199.40 1230.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,1184.70 C 1218.24,1191.00 1218.24,1199.40 1230.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,1184.70 C 1278.24,1191.00 1278.24,1199.40 1290.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,1184.70 C 1278.24,1191.00 1278.24,1199.40 1290.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,1184.70 C 1278.24,1191.00 1278.24,1199.40 1290.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,1184.70 C 1338.24,1191.00 1338.24,1199.40 1350.00,1205.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,1184.70 C 1338.24,1191.00 1338.24,1199.40 1350.00,1205.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,1184.70 C 1338.24,1191.00 1338.24,1199.40 1350.00,1205.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,1244.70 C 138.24,1251.00 138.24,1259.40 150.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,1244.70 C 138.24,1251.00 138.24,1259.40 150.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,1244.70 C 138.24,1251.00 138.24,1259.40 150.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,1244.70 C 198.24,1251.00 198.24,1259.40 210.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,1244.70 C 198.24,1251.00 198.24,1259.40 210.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,1244.70 C 198.24,1251.00 198.24,1259.40 210.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,1244.70 C 258.24,1251.00 258.24,1259.40 270.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,1244.70 C 258.24,1251.00 258.24,1259.40 270.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,1244.70 C 258.24,1251.00 258.24,1259.40 270.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,1244.70 C 318.24,1251.00 318.24,1259.40 330.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,1244.70 C 318.24,1251.00 318.24,1259.40 330.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,1244.70 C 318.24,1251.00 318.24,1259.40 330.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,1244.70 C 378.24,1251.00 378.24,1259.40 390.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,1244.70 C 378.24,1251.00 378.24,1259.40 390.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,1244.70 C 378.24,1251.00 378.24,1259.40 390.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,1244.70 C 438.24,1251.00 438.24,1259.40 450.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,1244.70 C 438.24,1251.00 438.24,1259.40 450.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,1244.70 C 438.24,1251.00 438.24,1259.40 450.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,1244.70 C 498.24,1251.00 498.24,1259.40 510.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,1244.70 C 498.24,1251.00 498.24,1259.40 510.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,1244.70 C 498.24,1251.00 498.24,1259.40 510.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,1244.70 C 558.24,1251.00 558.24,1259.40 570.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,1244.70 C 558.24,1251.00 558.24,1259.40 570.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,1244.70 C 558.24,1251.00 558.24,1259.40 570.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,1244.70 C 618.24,1251.00 618.24,1259.40 630.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,1244.70 C 618.24,1251.00 618.24,1259.40 630.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,1244.70 C 618.24,1251.00 618.24,1259.40 630.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,1244.70 C 678.24,1251.00 678.24,1259.40 690.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,1244.70 C 678.24,1251.00 678.24,1259.40 690.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,1244.70 C 678.24,1251.00 678.24,1259.40 690.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,1244.70 C 738.24,1251.00 738.24,1259.40 750.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,1244.70 C 738.24,1251.00 738.24,1259.40 750.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,1244.70 C 738.24,1251.00 738.24,1259.40 750.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,1244.70 C 798.24,1251.00 798.24,1259.40 810.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,1244.70 C 798.24,1251.00 798.24,1259.40 810.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,1244.70 C 798.24,1251.00 798.24,1259.40 810.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,1244.70 C 858.24,1251.00 858.24,1259.40 870.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,1244.70 C 858.24,1251.00 858.24,1259.40 870.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,1244.70 C 858.24,1251.00 858.24,1259.40 870.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,1244.70 C 918.24,1251.00 918.24,1259.40 930.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,1244.70 C 918.24,1251.00 918.24,1259.40 930.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,1244.70 C 918.24,1251.00 918.24,1259.40 930.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,1244.70 C 978.24,1251.00 978.24,1259.40 990.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,1244.70 C 978.24,1251.00 978.24,1259.40 990.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,1244.70 C 978.24,1251.00 978.24,1259.40 990.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,1244.70 C 1038.24,1251.00 1038.24,1259.40 1050.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,1244.70 C 1038.24,1251.00 1038.24,1259.40 1050.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,1244.70 C 1038.24,1251.00 1038.24,1259.40 1050.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,1244.70 C 1098.24,1251.00 1098.24,1259.40 1110.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,1244.70 C 1098.24,1251.00 1098.24,1259.40 1110.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,1244.70 C 1098.24,1251.00 1098.24,1259.40 1110.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,1244.70 C 1158.24,1251.00 1158.24,1259.40 1170.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,1244.70 C 1158.24,1251.00 1158.24,1259.40 1170.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,1244.70 C 1158.24,1251.00 1158.24,1259.40 1170.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,1244.70 C 1218.24,1251.00 1218.24,1259.40 1230.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,1244.70 C 1218.24,1251.00 1218.24,1259.40 1230.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,1244.70 C 1218.24,1251.00 1218.24,1259.40 1230.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,1244.70 C 1278.24,1251.00 1278.24,1259.40 1290.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,1244.70 C 1278.24,1251.00 1278.24,1259.40 1290.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,1244.70 C 1278.24,1251.00 1278.24,1259.40 1290.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,1244.70 C 1338.24,1251.00 1338.24,1259.40 1350.00,1265.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,1244.70 C 1338.24,1251.00 1338.24,1259.40 1350.00,1265.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,1244.70 C 1338.24,1251.00 1338.24,1259.40 1350.00,1265.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 150.00,1304.70 C 138.24,1311.00 138.24,1319.40 150.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 150.00,1304.70 C 138.24,1311.00 138.24,1319.40 150.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 150.00,1304.70 C 138.24,1311.00 138.24,1319.40 150.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 210.00,1304.70 C 198.24,1311.00 198.24,1319.40 210.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 210.00,1304.70 C 198.24,1311.00 198.24,1319.40 210.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 210.00,1304.70 C 198.24,1311.00 198.24,1319.40 210.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 270.00,1304.70 C 258.24,1311.00 258.24,1319.40 270.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 270.00,1304.70 C 258.24,1311.00 258.24,1319.40 270.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 270.00,1304.70 C 258.24,1311.00 258.24,1319.40 270.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 330.00,1304.70 C 318.24,1311.00 318.24,1319.40 330.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 330.00,1304.70 C 318.24,1311.00 318.24,1319.40 330.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 330.00,1304.70 C 318.24,1311.00 318.24,1319.40 330.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 390.00,1304.70 C 378.24,1311.00 378.24,1319.40 390.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 390.00,1304.70 C 378.24,1311.00 378.24,1319.40 390.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 390.00,1304.70 C 378.24,1311.00 378.24,1319.40 390.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 450.00,1304.70 C 438.24,1311.00 438.24,1319.40 450.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 450.00,1304.70 C 438.24,1311.00 438.24,1319.40 450.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 450.00,1304.70 C 438.24,1311.00 438.24,1319.40 450.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 510.00,1304.70 C 498.24,1311.00 498.24,1319.40 510.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 510.00,1304.70 C 498.24,1311.00 498.24,1319.40 510.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 510.00,1304.70 C 498.24,1311.00 498.24,1319.40 510.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 570.00,1304.70 C 558.24,1311.00 558.24,1319.40 570.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 570.00,1304.70 C 558.24,1311.00 558.24,1319.40 570.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 570.00,1304.70 C 558.24,1311.00 558.24,1319.40 570.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 630.00,1304.70 C 618.24,1311.00 618.24,1319.40 630.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 630.00,1304.70 C 618.24,1311.00 618.24,1319.40 630.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 630.00,1304.70 C 618.24,1311.00 618.24,1319.40 630.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 690.00,1304.70 C 678.24,1311.00 678.24,1319.40 690.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 690.00,1304.70 C 678.24,1311.00 678.24,1319.40 690.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 690.00,1304.70 C 678.24,1311.00 678.24,1319.40 690.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 750.00,1304.70 C 738.24,1311.00 738.24,1319.40 750.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 750.00,1304.70 C 738.24,1311.00 738.24,1319.40 750.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 750.00,1304.70 C 738.24,1311.00 738.24,1319.40 750.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 810.00,1304.70 C 798.24,1311.00 798.24,1319.40 810.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 810.00,1304.70 C 798.24,1311.00 798.24,1319.40 810.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 810.00,1304.70 C 798.24,1311.00 798.24,1319.40 810.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 870.00,1304.70 C 858.24,1311.00 858.24,1319.40 870.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 870.00,1304.70 C 858.24,1311.00 858.24,1319.40 870.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 870.00,1304.70 C 858.24,1311.00 858.24,1319.40 870.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 930.00,1304.70 C 918.24,1311.00 918.24,1319.40 930.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 930.00,1304.70 C 918.24,1311.00 918.24,1319.40 930.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 930.00,1304.70 C 918.24,1311.00 918.24,1319.40 930.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 990.00,1304.70 C 978.24,1311.00 978.24,1319.40 990.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 990.00,1304.70 C 978.24,1311.00 978.24,1319.40 990.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 990.00,1304.70 C 978.24,1311.00 978.24,1319.40 990.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1050.00,1304.70 C 1038.24,1311.00 1038.24,1319.40 1050.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1050.00,1304.70 C 1038.24,1311.00 1038.24,1319.40 1050.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1050.00,1304.70 C 1038.24,1311.00 1038.24,1319.40 1050.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1110.00,1304.70 C 1098.24,1311.00 1098.24,1319.40 1110.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1110.00,1304.70 C 1098.24,1311.00 1098.24,1319.40 1110.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1110.00,1304.70 C 1098.24,1311.00 1098.24,1319.40 1110.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1170.00,1304.70 C 1158.24,1311.00 1158.24,1319.40 1170.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1170.00,1304.70 C 1158.24,1311.00 1158.24,1319.40 1170.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1170.00,1304.70 C 1158.24,1311.00 1158.24,1319.40 1170.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1230.00,1304.70 C 1218.24,1311.00 1218.24,1319.40 1230.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1230.00,1304.70 C 1218.24,1311.00 1218.24,1319.40 1230.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1230.00,1304.70 C 1218.24,1311.00 1218.24,1319.40 1230.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1290.00,1304.70 C 1278.24,1311.00 1278.24,1319.40 1290.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1290.00,1304.70 C 1278.24,1311.00 1278.24,1319.40 1290.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1290.00,1304.70 C 1278.24,1311.00 1278.24,1319.40 1290.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /><path d="M 1350.00,1304.70 C 1338.24,1311.00 1338.24,1319.40 1350.00,1325.70" fill="none" stroke="#000000" stroke-linecap="round" stroke-linejoin="round" stroke-opacity="0.3" stroke-width="7.919999999999999" transform="translate(0.5,0.5)" /><path d="M 1350.00,1304.70 C 1338.24,1311.00 1338.24,1319.40 1350.00,1325.70" fill="none" filter="url(#emboss)" stroke="url(#ropegrad)" stroke-linecap="round" stroke-linejoin="round" stroke-width="6.6" /><path d="M 1350.00,1304.70 C 1338.24,1311.00 1338.24,1319.40 1350.00,1325.70" fill="none" filter="url(#glow)" opacity="0.7" stroke="#ffffff" stroke-linecap="round" stroke-linejoin="round" stroke-width="4.2" /></g><g><path d="M 121.50,150.00 A 28.50,28.50 0 0 1 150.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 178.50,150.00 A 28.50,28.50 0 0 1 150.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,150.00 A 28.50,28.50 0 0 1 210.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 238.50,150.00 A 28.50,28.50 0 0 1 210.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,121.50 A 28.50,28.50 0 0 1 298.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,178.50 A 28.50,28.50 0 0 1 241.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,150.00 A 28.50,28.50 0 0 1 330.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,150.00 A 28.50,28.50 0 0 1 330.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,150.00 A 28.50,28.50 0 0 1 390.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,150.00 A 28.50,28.50 0 0 1 390.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,178.50 A 28.50,28.50 0 0 1 421.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,121.50 A 28.50,28.50 0 0 1 478.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,178.50 A 28.50,28.50 0 0 1 481.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,121.50 A 28.50,28.50 0 0 1 538.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="150.0" fill="black" r="3.5999999999999996" /><path d="M 541.50,150.00 A 28.50,28.50 0 0 1 570.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,150.00 A 28.50,28.50 0 0 1 570.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="570.0" cy="150.0" fill="black" r="3.5999999999999996" /><path d="M 601.50,150.00 A 28.50,28.50 0 0 1 630.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,150.00 A 28.50,28.50 0 0 1 630.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,150.00 A 28.50,28.50 0 0 1 690.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,150.00 A 28.50,28.50 0 0 1 690.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,150.00 A 28.50,28.50 0 0 1 750.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 778.50,150.00 A 28.50,28.50 0 0 1 750.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,150.00 A 28.50,28.50 0 0 1 810.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,150.00 A 28.50,28.50 0 0 1 810.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,150.00 A 28.50,28.50 0 0 1 870.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,150.00 A 28.50,28.50 0 0 1 870.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,150.00 A 28.50,28.50 0 0 1 930.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,150.00 A 28.50,28.50 0 0 1 930.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 961.50,150.00 A 28.50,28.50 0 0 1 990.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1018.50,150.00 A 28.50,28.50 0 0 1 990.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,150.00 A 28.50,28.50 0 0 1 1050.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,150.00 A 28.50,28.50 0 0 1 1050.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,121.50 A 28.50,28.50 0 0 1 1138.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,178.50 A 28.50,28.50 0 0 1 1081.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1110.0" cy="150.0" fill="black" r="3.5999999999999996" /><path d="M 1170.00,178.50 A 28.50,28.50 0 0 1 1141.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,121.50 A 28.50,28.50 0 0 1 1198.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,178.50 A 28.50,28.50 0 0 1 1201.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,121.50 A 28.50,28.50 0 0 1 1258.50,150.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,150.00 A 28.50,28.50 0 0 1 1290.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,150.00 A 28.50,28.50 0 0 1 1290.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1290.0" cy="150.0" fill="black" r="3.5999999999999996" /><path d="M 1321.50,150.00 A 28.50,28.50 0 0 1 1350.00,121.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,150.00 A 28.50,28.50 0 0 1 1350.00,178.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1350.0" cy="150.0" fill="black" r="3.5999999999999996" /><path d="M 178.50,210.00 A 28.50,28.50 0 0 1 150.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 121.50,210.00 A 28.50,28.50 0 0 1 150.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 210.00,238.50 A 28.50,28.50 0 0 1 181.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,181.50 A 28.50,28.50 0 0 1 238.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 298.50,210.00 A 28.50,28.50 0 0 1 270.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 241.50,210.00 A 28.50,28.50 0 0 1 270.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="270.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 330.00,181.50 A 28.50,28.50 0 0 1 358.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,238.50 A 28.50,28.50 0 0 1 301.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="330.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 361.50,210.00 A 28.50,28.50 0 0 1 390.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,210.00 A 28.50,28.50 0 0 1 390.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,210.00 A 28.50,28.50 0 0 1 450.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,210.00 A 28.50,28.50 0 0 1 450.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,238.50 A 28.50,28.50 0 0 1 481.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,181.50 A 28.50,28.50 0 0 1 538.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 570.00,181.50 A 28.50,28.50 0 0 1 598.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,238.50 A 28.50,28.50 0 0 1 541.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,210.00 A 28.50,28.50 0 0 1 630.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,210.00 A 28.50,28.50 0 0 1 630.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="630.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 718.50,210.00 A 28.50,28.50 0 0 1 690.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,210.00 A 28.50,28.50 0 0 1 690.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="690.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 778.50,210.00 A 28.50,28.50 0 0 1 750.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,210.00 A 28.50,28.50 0 0 1 750.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,181.50 A 28.50,28.50 0 0 1 838.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,238.50 A 28.50,28.50 0 0 1 781.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="810.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 841.50,210.00 A 28.50,28.50 0 0 1 870.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,210.00 A 28.50,28.50 0 0 1 870.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 930.00,181.50 A 28.50,28.50 0 0 1 958.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,238.50 A 28.50,28.50 0 0 1 901.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,181.50 A 28.50,28.50 0 0 1 1018.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,238.50 A 28.50,28.50 0 0 1 961.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,210.00 A 28.50,28.50 0 0 1 1050.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,210.00 A 28.50,28.50 0 0 1 1050.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,210.00 A 28.50,28.50 0 0 1 1110.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1138.50,210.00 A 28.50,28.50 0 0 1 1110.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1110.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 1198.50,210.00 A 28.50,28.50 0 0 1 1170.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1141.50,210.00 A 28.50,28.50 0 0 1 1170.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,210.00 A 28.50,28.50 0 0 1 1230.00,238.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1201.50,210.00 A 28.50,28.50 0 0 1 1230.00,181.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,181.50 A 28.50,28.50 0 0 1 1318.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,238.50 A 28.50,28.50 0 0 1 1261.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1290.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 1350.00,181.50 A 28.50,28.50 0 0 1 1378.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,238.50 A 28.50,28.50 0 0 1 1321.50,210.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1350.0" cy="210.0" fill="black" r="3.5999999999999996" /><path d="M 150.00,298.50 A 28.50,28.50 0 0 1 121.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,241.50 A 28.50,28.50 0 0 1 178.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,298.50 A 28.50,28.50 0 0 1 181.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,241.50 A 28.50,28.50 0 0 1 238.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="210.0" cy="270.0" fill="black" r="3.5999999999999996" /><path d="M 270.00,241.50 A 28.50,28.50 0 0 1 298.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,298.50 A 28.50,28.50 0 0 1 241.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,270.00 A 28.50,28.50 0 0 1 330.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,270.00 A 28.50,28.50 0 0 1 330.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="330.0" cy="270.0" fill="black" r="3.5999999999999996" /><path d="M 390.00,298.50 A 28.50,28.50 0 0 1 361.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,241.50 A 28.50,28.50 0 0 1 418.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,241.50 A 28.50,28.50 0 0 1 478.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,298.50 A 28.50,28.50 0 0 1 421.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="450.0" cy="270.0" fill="black" r="3.5999999999999996" /><path d="M 481.50,270.00 A 28.50,28.50 0 0 1 510.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 538.50,270.00 A 28.50,28.50 0 0 1 510.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="270.0" fill="black" r="3.5999999999999996" /><path d="M 541.50,270.00 A 28.50,28.50 0 0 1 570.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,270.00 A 28.50,28.50 0 0 1 570.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,270.00 A 28.50,28.50 0 0 1 630.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,270.00 A 28.50,28.50 0 0 1 630.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,298.50 A 28.50,28.50 0 0 1 661.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,241.50 A 28.50,28.50 0 0 1 718.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="690.0" cy="270.0" fill="black" r="3.5999999999999996" /><path d="M 750.00,241.50 A 28.50,28.50 0 0 1 778.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,298.50 A 28.50,28.50 0 0 1 721.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,270.00 A 28.50,28.50 0 0 1 810.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,270.00 A 28.50,28.50 0 0 1 810.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="810.0" cy="270.0" fill="black" r="3.5999999999999996" /><path d="M 898.50,270.00 A 28.50,28.50 0 0 1 870.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,270.00 A 28.50,28.50 0 0 1 870.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,270.00 A 28.50,28.50 0 0 1 930.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,270.00 A 28.50,28.50 0 0 1 930.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="270.0" fill="black" r="3.5999999999999996" /><path d="M 990.00,241.50 A 28.50,28.50 0 0 1 1018.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,298.50 A 28.50,28.50 0 0 1 961.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="990.0" cy="270.0" fill="black" r="3.5999999999999996" /><path d="M 1078.50,270.00 A 28.50,28.50 0 0 1 1050.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,270.00 A 28.50,28.50 0 0 1 1050.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,298.50 A 28.50,28.50 0 0 1 1081.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,241.50 A 28.50,28.50 0 0 1 1138.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,298.50 A 28.50,28.50 0 0 1 1141.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,241.50 A 28.50,28.50 0 0 1 1198.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1170.0" cy="270.0" fill="black" r="3.5999999999999996" /><path d="M 1230.00,241.50 A 28.50,28.50 0 0 1 1258.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,298.50 A 28.50,28.50 0 0 1 1201.50,270.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,270.00 A 28.50,28.50 0 0 1 1290.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,270.00 A 28.50,28.50 0 0 1 1290.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,270.00 A 28.50,28.50 0 0 1 1350.00,298.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,270.00 A 28.50,28.50 0 0 1 1350.00,241.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 121.50,330.00 A 28.50,28.50 0 0 1 150.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 178.50,330.00 A 28.50,28.50 0 0 1 150.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,301.50 A 28.50,28.50 0 0 1 238.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,358.50 A 28.50,28.50 0 0 1 181.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="210.0" cy="330.0" fill="black" r="3.5999999999999996" /><path d="M 298.50,330.00 A 28.50,28.50 0 0 1 270.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 241.50,330.00 A 28.50,28.50 0 0 1 270.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,358.50 A 28.50,28.50 0 0 1 301.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,301.50 A 28.50,28.50 0 0 1 358.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,358.50 A 28.50,28.50 0 0 1 361.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,301.50 A 28.50,28.50 0 0 1 418.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,330.00 A 28.50,28.50 0 0 1 450.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,330.00 A 28.50,28.50 0 0 1 450.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="450.0" cy="330.0" fill="black" r="3.5999999999999996" /><path d="M 481.50,330.00 A 28.50,28.50 0 0 1 510.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 538.50,330.00 A 28.50,28.50 0 0 1 510.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="330.0" fill="black" r="3.5999999999999996" /><path d="M 598.50,330.00 A 28.50,28.50 0 0 1 570.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,330.00 A 28.50,28.50 0 0 1 570.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,330.00 A 28.50,28.50 0 0 1 630.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,330.00 A 28.50,28.50 0 0 1 630.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,301.50 A 28.50,28.50 0 0 1 718.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,358.50 A 28.50,28.50 0 0 1 661.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="690.0" cy="330.0" fill="black" r="3.5999999999999996" /><path d="M 750.00,301.50 A 28.50,28.50 0 0 1 778.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,358.50 A 28.50,28.50 0 0 1 721.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="750.0" cy="330.0" fill="black" r="3.5999999999999996" /><path d="M 838.50,330.00 A 28.50,28.50 0 0 1 810.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,330.00 A 28.50,28.50 0 0 1 810.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,358.50 A 28.50,28.50 0 0 1 841.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,301.50 A 28.50,28.50 0 0 1 898.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,330.00 A 28.50,28.50 0 0 1 930.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,330.00 A 28.50,28.50 0 0 1 930.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="330.0" fill="black" r="3.5999999999999996" /><path d="M 1018.50,330.00 A 28.50,28.50 0 0 1 990.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 961.50,330.00 A 28.50,28.50 0 0 1 990.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,330.00 A 28.50,28.50 0 0 1 1050.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,330.00 A 28.50,28.50 0 0 1 1050.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,330.00 A 28.50,28.50 0 0 1 1110.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1138.50,330.00 A 28.50,28.50 0 0 1 1110.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,301.50 A 28.50,28.50 0 0 1 1198.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,358.50 A 28.50,28.50 0 0 1 1141.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1170.0" cy="330.0" fill="black" r="3.5999999999999996" /><path d="M 1201.50,330.00 A 28.50,28.50 0 0 1 1230.00,301.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,330.00 A 28.50,28.50 0 0 1 1230.00,358.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1230.0" cy="330.0" fill="black" r="3.5999999999999996" /><path d="M 1290.00,301.50 A 28.50,28.50 0 0 1 1318.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,358.50 A 28.50,28.50 0 0 1 1261.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,358.50 A 28.50,28.50 0 0 1 1321.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,301.50 A 28.50,28.50 0 0 1 1378.50,330.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1350.0" cy="330.0" fill="black" r="3.5999999999999996" /><path d="M 150.00,361.50 A 28.50,28.50 0 0 1 178.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,418.50 A 28.50,28.50 0 0 1 121.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="390.0" fill="black" r="3.5999999999999996" /><path d="M 238.50,390.00 A 28.50,28.50 0 0 1 210.00,418.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,390.00 A 28.50,28.50 0 0 1 210.00,361.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 298.50,390.00 A 28.50,28.50 0 0 1 270.00,418.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 241.50,390.00 A 28.50,28.50 0 0 1 270.00,361.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,390.00 A 28.50,28.50 0 0 1 330.00,361.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,390.00 A 28.50,28.50 0 0 1 330.00,418.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,361.50 A 28.50,28.50 0 0 1 418.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,418.50 A 28.50,28.50 0 0 1 361.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="390.0" cy="390.0" fill="black" r="3.5999999999999996" /><path d="M 450.00,361.50 A 28.50,28.50 0 0 1 478.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,418.50 A 28.50,28.50 0 0 1 421.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,361.50 A 28.50,28.50 0 0 1 538.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,418.50 A 28.50,28.50 0 0 1 481.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,418.50 A 28.50,28.50 0 0 1 541.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,361.50 A 28.50,28.50 0 0 1 598.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,390.00 A 28.50,28.50 0 0 1 630.00,418.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,390.00 A 28.50,28.50 0 0 1 630.00,361.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="630.0" cy="390.0" fill="black" r="3.5999999999999996" /><path d="M 661.50,390.00 A 28.50,28.50 0 0 1 690.00,361.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,390.00 A 28.50,28.50 0 0 1 690.00,418.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="690.0" cy="390.0" fill="black" r="3.5999999999999996" /><path d="M 750.00,418.50 A 28.50,28.50 0 0 1 721.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,361.50 A 28.50,28.50 0 0 1 778.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,418.50 A 28.50,28.50 0 0 1 781.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,361.50 A 28.50,28.50 0 0 1 838.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="810.0" cy="390.0" fill="black" r="3.5999999999999996" /><path d="M 870.00,361.50 A 28.50,28.50 0 0 1 898.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,418.50 A 28.50,28.50 0 0 1 841.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="390.0" fill="black" r="3.5999999999999996" /><path d="M 901.50,390.00 A 28.50,28.50 0 0 1 930.00,361.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,390.00 A 28.50,28.50 0 0 1 930.00,418.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="390.0" fill="black" r="3.5999999999999996" /><path d="M 990.00,361.50 A 28.50,28.50 0 0 1 1018.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,418.50 A 28.50,28.50 0 0 1 961.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1050.00,361.50 A 28.50,28.50 0 0 1 1078.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1050.00,418.50 A 28.50,28.50 0 0 1 1021.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,390.00 A 28.50,28.50 0 0 1 1110.00,361.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1138.50,390.00 A 28.50,28.50 0 0 1 1110.00,418.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1141.50,390.00 A 28.50,28.50 0 0 1 1170.00,361.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,390.00 A 28.50,28.50 0 0 1 1170.00,418.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1170.0" cy="390.0" fill="black" r="3.5999999999999996" /><path d="M 1230.00,418.50 A 28.50,28.50 0 0 1 1201.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,361.50 A 28.50,28.50 0 0 1 1258.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,418.50 A 28.50,28.50 0 0 1 1261.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,361.50 A 28.50,28.50 0 0 1 1318.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,361.50 A 28.50,28.50 0 0 1 1378.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,418.50 A 28.50,28.50 0 0 1 1321.50,390.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1350.0" cy="390.0" fill="black" r="3.5999999999999996" /><path d="M 150.00,421.50 A 28.50,28.50 0 0 1 178.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,478.50 A 28.50,28.50 0 0 1 121.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 238.50,450.00 A 28.50,28.50 0 0 1 210.00,478.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,450.00 A 28.50,28.50 0 0 1 210.00,421.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,421.50 A 28.50,28.50 0 0 1 298.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,478.50 A 28.50,28.50 0 0 1 241.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,450.00 A 28.50,28.50 0 0 1 330.00,421.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,450.00 A 28.50,28.50 0 0 1 330.00,478.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,450.00 A 28.50,28.50 0 0 1 390.00,421.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,450.00 A 28.50,28.50 0 0 1 390.00,478.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="390.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 450.00,478.50 A 28.50,28.50 0 0 1 421.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,421.50 A 28.50,28.50 0 0 1 478.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,478.50 A 28.50,28.50 0 0 1 481.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,421.50 A 28.50,28.50 0 0 1 538.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 570.00,421.50 A 28.50,28.50 0 0 1 598.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,478.50 A 28.50,28.50 0 0 1 541.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="570.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 601.50,450.00 A 28.50,28.50 0 0 1 630.00,421.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,450.00 A 28.50,28.50 0 0 1 630.00,478.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="630.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 690.00,421.50 A 28.50,28.50 0 0 1 718.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,478.50 A 28.50,28.50 0 0 1 661.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,478.50 A 28.50,28.50 0 0 1 721.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,421.50 A 28.50,28.50 0 0 1 778.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,421.50 A 28.50,28.50 0 0 1 838.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,478.50 A 28.50,28.50 0 0 1 781.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="810.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 841.50,450.00 A 28.50,28.50 0 0 1 870.00,421.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,450.00 A 28.50,28.50 0 0 1 870.00,478.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 958.50,450.00 A 28.50,28.50 0 0 1 930.00,478.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,450.00 A 28.50,28.50 0 0 1 930.00,421.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 990.00,421.50 A 28.50,28.50 0 0 1 1018.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,478.50 A 28.50,28.50 0 0 1 961.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="990.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 1050.00,421.50 A 28.50,28.50 0 0 1 1078.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1050.00,478.50 A 28.50,28.50 0 0 1 1021.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1050.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 1110.00,421.50 A 28.50,28.50 0 0 1 1138.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,478.50 A 28.50,28.50 0 0 1 1081.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1110.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 1198.50,450.00 A 28.50,28.50 0 0 1 1170.00,478.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1141.50,450.00 A 28.50,28.50 0 0 1 1170.00,421.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,478.50 A 28.50,28.50 0 0 1 1201.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,421.50 A 28.50,28.50 0 0 1 1258.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1230.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 1290.00,421.50 A 28.50,28.50 0 0 1 1318.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,478.50 A 28.50,28.50 0 0 1 1261.50,450.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1290.0" cy="450.0" fill="black" r="3.5999999999999996" /><path d="M 1321.50,450.00 A 28.50,28.50 0 0 1 1350.00,421.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,450.00 A 28.50,28.50 0 0 1 1350.00,478.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 178.50,510.00 A 28.50,28.50 0 0 1 150.00,538.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 121.50,510.00 A 28.50,28.50 0 0 1 150.00,481.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,510.00 A 28.50,28.50 0 0 1 210.00,481.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 238.50,510.00 A 28.50,28.50 0 0 1 210.00,538.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,481.50 A 28.50,28.50 0 0 1 298.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,538.50 A 28.50,28.50 0 0 1 241.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="270.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 301.50,510.00 A 28.50,28.50 0 0 1 330.00,481.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,510.00 A 28.50,28.50 0 0 1 330.00,538.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="330.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 390.00,481.50 A 28.50,28.50 0 0 1 418.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,538.50 A 28.50,28.50 0 0 1 361.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,538.50 A 28.50,28.50 0 0 1 421.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,481.50 A 28.50,28.50 0 0 1 478.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="450.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 510.00,481.50 A 28.50,28.50 0 0 1 538.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,538.50 A 28.50,28.50 0 0 1 481.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 598.50,510.00 A 28.50,28.50 0 0 1 570.00,538.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,510.00 A 28.50,28.50 0 0 1 570.00,481.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="570.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 630.00,538.50 A 28.50,28.50 0 0 1 601.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,481.50 A 28.50,28.50 0 0 1 658.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,538.50 A 28.50,28.50 0 0 1 661.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,481.50 A 28.50,28.50 0 0 1 718.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,481.50 A 28.50,28.50 0 0 1 778.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,538.50 A 28.50,28.50 0 0 1 721.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="750.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 810.00,481.50 A 28.50,28.50 0 0 1 838.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,538.50 A 28.50,28.50 0 0 1 781.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,538.50 A 28.50,28.50 0 0 1 841.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,481.50 A 28.50,28.50 0 0 1 898.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,538.50 A 28.50,28.50 0 0 1 901.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,481.50 A 28.50,28.50 0 0 1 958.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,538.50 A 28.50,28.50 0 0 1 961.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,481.50 A 28.50,28.50 0 0 1 1018.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="990.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 1021.50,510.00 A 28.50,28.50 0 0 1 1050.00,481.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,510.00 A 28.50,28.50 0 0 1 1050.00,538.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1050.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 1110.00,538.50 A 28.50,28.50 0 0 1 1081.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,481.50 A 28.50,28.50 0 0 1 1138.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,538.50 A 28.50,28.50 0 0 1 1141.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,481.50 A 28.50,28.50 0 0 1 1198.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1170.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 1230.00,481.50 A 28.50,28.50 0 0 1 1258.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,538.50 A 28.50,28.50 0 0 1 1201.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1230.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 1261.50,510.00 A 28.50,28.50 0 0 1 1290.00,481.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,510.00 A 28.50,28.50 0 0 1 1290.00,538.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1290.0" cy="510.0" fill="black" r="3.5999999999999996" /><path d="M 1350.00,481.50 A 28.50,28.50 0 0 1 1378.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,538.50 A 28.50,28.50 0 0 1 1321.50,510.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,598.50 A 28.50,28.50 0 0 1 121.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,541.50 A 28.50,28.50 0 0 1 178.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 210.00,541.50 A 28.50,28.50 0 0 1 238.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,598.50 A 28.50,28.50 0 0 1 181.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="210.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 241.50,570.00 A 28.50,28.50 0 0 1 270.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 298.50,570.00 A 28.50,28.50 0 0 1 270.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="270.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 358.50,570.00 A 28.50,28.50 0 0 1 330.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,570.00 A 28.50,28.50 0 0 1 330.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="330.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 390.00,541.50 A 28.50,28.50 0 0 1 418.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,598.50 A 28.50,28.50 0 0 1 361.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="390.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 450.00,541.50 A 28.50,28.50 0 0 1 478.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,598.50 A 28.50,28.50 0 0 1 421.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="450.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 510.00,541.50 A 28.50,28.50 0 0 1 538.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,598.50 A 28.50,28.50 0 0 1 481.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 598.50,570.00 A 28.50,28.50 0 0 1 570.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,570.00 A 28.50,28.50 0 0 1 570.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,598.50 A 28.50,28.50 0 0 1 601.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,541.50 A 28.50,28.50 0 0 1 658.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="630.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 690.00,541.50 A 28.50,28.50 0 0 1 718.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,598.50 A 28.50,28.50 0 0 1 661.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="690.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 778.50,570.00 A 28.50,28.50 0 0 1 750.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,570.00 A 28.50,28.50 0 0 1 750.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="750.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 838.50,570.00 A 28.50,28.50 0 0 1 810.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,570.00 A 28.50,28.50 0 0 1 810.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="810.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 870.00,541.50 A 28.50,28.50 0 0 1 898.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,598.50 A 28.50,28.50 0 0 1 841.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 930.00,541.50 A 28.50,28.50 0 0 1 958.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,598.50 A 28.50,28.50 0 0 1 901.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 961.50,570.00 A 28.50,28.50 0 0 1 990.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1018.50,570.00 A 28.50,28.50 0 0 1 990.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,570.00 A 28.50,28.50 0 0 1 1050.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,570.00 A 28.50,28.50 0 0 1 1050.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,598.50 A 28.50,28.50 0 0 1 1081.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,541.50 A 28.50,28.50 0 0 1 1138.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1110.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 1170.00,541.50 A 28.50,28.50 0 0 1 1198.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,598.50 A 28.50,28.50 0 0 1 1141.50,570.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1170.0" cy="570.0" fill="black" r="3.5999999999999996" /><path d="M 1201.50,570.00 A 28.50,28.50 0 0 1 1230.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,570.00 A 28.50,28.50 0 0 1 1230.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,570.00 A 28.50,28.50 0 0 1 1290.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,570.00 A 28.50,28.50 0 0 1 1290.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,570.00 A 28.50,28.50 0 0 1 1350.00,541.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,570.00 A 28.50,28.50 0 0 1 1350.00,598.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,601.50 A 28.50,28.50 0 0 1 178.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,658.50 A 28.50,28.50 0 0 1 121.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="630.0" fill="black" r="3.5999999999999996" /><path d="M 238.50,630.00 A 28.50,28.50 0 0 1 210.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,630.00 A 28.50,28.50 0 0 1 210.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="210.0" cy="630.0" fill="black" r="3.5999999999999996" /><path d="M 270.00,658.50 A 28.50,28.50 0 0 1 241.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,601.50 A 28.50,28.50 0 0 1 298.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,658.50 A 28.50,28.50 0 0 1 301.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,601.50 A 28.50,28.50 0 0 1 358.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,601.50 A 28.50,28.50 0 0 1 418.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,658.50 A 28.50,28.50 0 0 1 361.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,630.00 A 28.50,28.50 0 0 1 450.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,630.00 A 28.50,28.50 0 0 1 450.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="450.0" cy="630.0" fill="black" r="3.5999999999999996" /><path d="M 538.50,630.00 A 28.50,28.50 0 0 1 510.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 481.50,630.00 A 28.50,28.50 0 0 1 510.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="630.0" fill="black" r="3.5999999999999996" /><path d="M 570.00,658.50 A 28.50,28.50 0 0 1 541.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,601.50 A 28.50,28.50 0 0 1 598.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,601.50 A 28.50,28.50 0 0 1 658.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,658.50 A 28.50,28.50 0 0 1 601.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="630.0" cy="630.0" fill="black" r="3.5999999999999996" /><path d="M 718.50,630.00 A 28.50,28.50 0 0 1 690.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,630.00 A 28.50,28.50 0 0 1 690.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="690.0" cy="630.0" fill="black" r="3.5999999999999996" /><path d="M 778.50,630.00 A 28.50,28.50 0 0 1 750.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,630.00 A 28.50,28.50 0 0 1 750.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,658.50 A 28.50,28.50 0 0 1 781.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,601.50 A 28.50,28.50 0 0 1 838.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,630.00 A 28.50,28.50 0 0 1 870.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,630.00 A 28.50,28.50 0 0 1 870.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="630.0" fill="black" r="3.5999999999999996" /><path d="M 958.50,630.00 A 28.50,28.50 0 0 1 930.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,630.00 A 28.50,28.50 0 0 1 930.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="630.0" fill="black" r="3.5999999999999996" /><path d="M 990.00,658.50 A 28.50,28.50 0 0 1 961.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,601.50 A 28.50,28.50 0 0 1 1018.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1050.00,658.50 A 28.50,28.50 0 0 1 1021.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1050.00,601.50 A 28.50,28.50 0 0 1 1078.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,630.00 A 28.50,28.50 0 0 1 1110.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1138.50,630.00 A 28.50,28.50 0 0 1 1110.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1110.0" cy="630.0" fill="black" r="3.5999999999999996" /><path d="M 1141.50,630.00 A 28.50,28.50 0 0 1 1170.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,630.00 A 28.50,28.50 0 0 1 1170.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1201.50,630.00 A 28.50,28.50 0 0 1 1230.00,601.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,630.00 A 28.50,28.50 0 0 1 1230.00,658.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,658.50 A 28.50,28.50 0 0 1 1261.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,601.50 A 28.50,28.50 0 0 1 1318.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,601.50 A 28.50,28.50 0 0 1 1378.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,658.50 A 28.50,28.50 0 0 1 1321.50,630.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 178.50,690.00 A 28.50,28.50 0 0 1 150.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 121.50,690.00 A 28.50,28.50 0 0 1 150.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 238.50,690.00 A 28.50,28.50 0 0 1 210.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,690.00 A 28.50,28.50 0 0 1 210.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="210.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 270.00,661.50 A 28.50,28.50 0 0 1 298.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,718.50 A 28.50,28.50 0 0 1 241.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="270.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 330.00,661.50 A 28.50,28.50 0 0 1 358.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,718.50 A 28.50,28.50 0 0 1 301.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="330.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 418.50,690.00 A 28.50,28.50 0 0 1 390.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,690.00 A 28.50,28.50 0 0 1 390.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="390.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 478.50,690.00 A 28.50,28.50 0 0 1 450.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,690.00 A 28.50,28.50 0 0 1 450.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,718.50 A 28.50,28.50 0 0 1 481.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,661.50 A 28.50,28.50 0 0 1 538.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,661.50 A 28.50,28.50 0 0 1 598.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,718.50 A 28.50,28.50 0 0 1 541.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,690.00 A 28.50,28.50 0 0 1 630.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,690.00 A 28.50,28.50 0 0 1 630.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,690.00 A 28.50,28.50 0 0 1 690.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,690.00 A 28.50,28.50 0 0 1 690.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,690.00 A 28.50,28.50 0 0 1 750.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 778.50,690.00 A 28.50,28.50 0 0 1 750.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,661.50 A 28.50,28.50 0 0 1 838.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 810.00,718.50 A 28.50,28.50 0 0 1 781.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="810.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 898.50,690.00 A 28.50,28.50 0 0 1 870.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,690.00 A 28.50,28.50 0 0 1 870.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 930.00,718.50 A 28.50,28.50 0 0 1 901.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,661.50 A 28.50,28.50 0 0 1 958.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,718.50 A 28.50,28.50 0 0 1 961.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,661.50 A 28.50,28.50 0 0 1 1018.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,690.00 A 28.50,28.50 0 0 1 1050.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,690.00 A 28.50,28.50 0 0 1 1050.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1050.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 1138.50,690.00 A 28.50,28.50 0 0 1 1110.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,690.00 A 28.50,28.50 0 0 1 1110.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1110.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 1170.00,718.50 A 28.50,28.50 0 0 1 1141.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,661.50 A 28.50,28.50 0 0 1 1198.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,718.50 A 28.50,28.50 0 0 1 1201.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,661.50 A 28.50,28.50 0 0 1 1258.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1230.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 1290.00,661.50 A 28.50,28.50 0 0 1 1318.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,718.50 A 28.50,28.50 0 0 1 1261.50,690.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1290.0" cy="690.0" fill="black" r="3.5999999999999996" /><path d="M 1378.50,690.00 A 28.50,28.50 0 0 1 1350.00,718.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,690.00 A 28.50,28.50 0 0 1 1350.00,661.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,721.50 A 28.50,28.50 0 0 1 178.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,778.50 A 28.50,28.50 0 0 1 121.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,778.50 A 28.50,28.50 0 0 1 181.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,721.50 A 28.50,28.50 0 0 1 238.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,778.50 A 28.50,28.50 0 0 1 241.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,721.50 A 28.50,28.50 0 0 1 298.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="270.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 358.50,750.00 A 28.50,28.50 0 0 1 330.00,778.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,750.00 A 28.50,28.50 0 0 1 330.00,721.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="330.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 418.50,750.00 A 28.50,28.50 0 0 1 390.00,778.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,750.00 A 28.50,28.50 0 0 1 390.00,721.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="390.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 450.00,721.50 A 28.50,28.50 0 0 1 478.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,778.50 A 28.50,28.50 0 0 1 421.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,721.50 A 28.50,28.50 0 0 1 538.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,778.50 A 28.50,28.50 0 0 1 481.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 541.50,750.00 A 28.50,28.50 0 0 1 570.00,721.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,750.00 A 28.50,28.50 0 0 1 570.00,778.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="570.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 630.00,721.50 A 28.50,28.50 0 0 1 658.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,778.50 A 28.50,28.50 0 0 1 601.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,778.50 A 28.50,28.50 0 0 1 661.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,721.50 A 28.50,28.50 0 0 1 718.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 778.50,750.00 A 28.50,28.50 0 0 1 750.00,778.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,750.00 A 28.50,28.50 0 0 1 750.00,721.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="750.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 838.50,750.00 A 28.50,28.50 0 0 1 810.00,778.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,750.00 A 28.50,28.50 0 0 1 810.00,721.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="810.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 870.00,778.50 A 28.50,28.50 0 0 1 841.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,721.50 A 28.50,28.50 0 0 1 898.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,778.50 A 28.50,28.50 0 0 1 901.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,721.50 A 28.50,28.50 0 0 1 958.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 990.00,721.50 A 28.50,28.50 0 0 1 1018.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,778.50 A 28.50,28.50 0 0 1 961.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="990.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 1078.50,750.00 A 28.50,28.50 0 0 1 1050.00,778.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,750.00 A 28.50,28.50 0 0 1 1050.00,721.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,721.50 A 28.50,28.50 0 0 1 1138.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,778.50 A 28.50,28.50 0 0 1 1081.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,778.50 A 28.50,28.50 0 0 1 1141.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,721.50 A 28.50,28.50 0 0 1 1198.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,721.50 A 28.50,28.50 0 0 1 1258.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,778.50 A 28.50,28.50 0 0 1 1201.50,750.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,750.00 A 28.50,28.50 0 0 1 1290.00,778.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,750.00 A 28.50,28.50 0 0 1 1290.00,721.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1290.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 1378.50,750.00 A 28.50,28.50 0 0 1 1350.00,778.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,750.00 A 28.50,28.50 0 0 1 1350.00,721.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1350.0" cy="750.0" fill="black" r="3.5999999999999996" /><path d="M 150.00,838.50 A 28.50,28.50 0 0 1 121.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,781.50 A 28.50,28.50 0 0 1 178.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,781.50 A 28.50,28.50 0 0 1 238.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,838.50 A 28.50,28.50 0 0 1 181.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="210.0" cy="810.0" fill="black" r="3.5999999999999996" /><path d="M 270.00,781.50 A 28.50,28.50 0 0 1 298.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,838.50 A 28.50,28.50 0 0 1 241.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,838.50 A 28.50,28.50 0 0 1 301.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,781.50 A 28.50,28.50 0 0 1 358.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,781.50 A 28.50,28.50 0 0 1 418.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,838.50 A 28.50,28.50 0 0 1 361.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="390.0" cy="810.0" fill="black" r="3.5999999999999996" /><path d="M 421.50,810.00 A 28.50,28.50 0 0 1 450.00,781.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,810.00 A 28.50,28.50 0 0 1 450.00,838.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="450.0" cy="810.0" fill="black" r="3.5999999999999996" /><path d="M 481.50,810.00 A 28.50,28.50 0 0 1 510.00,781.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 538.50,810.00 A 28.50,28.50 0 0 1 510.00,838.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,838.50 A 28.50,28.50 0 0 1 541.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,781.50 A 28.50,28.50 0 0 1 598.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,810.00 A 28.50,28.50 0 0 1 630.00,838.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,810.00 A 28.50,28.50 0 0 1 630.00,781.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,781.50 A 28.50,28.50 0 0 1 718.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,838.50 A 28.50,28.50 0 0 1 661.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="690.0" cy="810.0" fill="black" r="3.5999999999999996" /><path d="M 778.50,810.00 A 28.50,28.50 0 0 1 750.00,838.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,810.00 A 28.50,28.50 0 0 1 750.00,781.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,810.00 A 28.50,28.50 0 0 1 810.00,838.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,810.00 A 28.50,28.50 0 0 1 810.00,781.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,781.50 A 28.50,28.50 0 0 1 898.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,838.50 A 28.50,28.50 0 0 1 841.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="810.0" fill="black" r="3.5999999999999996" /><path d="M 901.50,810.00 A 28.50,28.50 0 0 1 930.00,781.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,810.00 A 28.50,28.50 0 0 1 930.00,838.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="810.0" fill="black" r="3.5999999999999996" /><path d="M 961.50,810.00 A 28.50,28.50 0 0 1 990.00,781.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1018.50,810.00 A 28.50,28.50 0 0 1 990.00,838.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1050.00,838.50 A 28.50,28.50 0 0 1 1021.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1050.00,781.50 A 28.50,28.50 0 0 1 1078.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,781.50 A 28.50,28.50 0 0 1 1138.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,838.50 A 28.50,28.50 0 0 1 1081.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1110.0" cy="810.0" fill="black" r="3.5999999999999996" /><path d="M 1170.00,781.50 A 28.50,28.50 0 0 1 1198.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,838.50 A 28.50,28.50 0 0 1 1141.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1170.0" cy="810.0" fill="black" r="3.5999999999999996" /><path d="M 1258.50,810.00 A 28.50,28.50 0 0 1 1230.00,838.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1201.50,810.00 A 28.50,28.50 0 0 1 1230.00,781.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,810.00 A 28.50,28.50 0 0 1 1290.00,838.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,810.00 A 28.50,28.50 0 0 1 1290.00,781.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,838.50 A 28.50,28.50 0 0 1 1321.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,781.50 A 28.50,28.50 0 0 1 1378.50,810.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,841.50 A 28.50,28.50 0 0 1 178.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,898.50 A 28.50,28.50 0 0 1 121.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="870.0" fill="black" r="3.5999999999999996" /><path d="M 181.50,870.00 A 28.50,28.50 0 0 1 210.00,841.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 238.50,870.00 A 28.50,28.50 0 0 1 210.00,898.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,898.50 A 28.50,28.50 0 0 1 241.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,841.50 A 28.50,28.50 0 0 1 298.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,841.50 A 28.50,28.50 0 0 1 358.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,898.50 A 28.50,28.50 0 0 1 301.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,870.00 A 28.50,28.50 0 0 1 390.00,841.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,870.00 A 28.50,28.50 0 0 1 390.00,898.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="390.0" cy="870.0" fill="black" r="3.5999999999999996" /><path d="M 478.50,870.00 A 28.50,28.50 0 0 1 450.00,898.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,870.00 A 28.50,28.50 0 0 1 450.00,841.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,898.50 A 28.50,28.50 0 0 1 481.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,841.50 A 28.50,28.50 0 0 1 538.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,841.50 A 28.50,28.50 0 0 1 598.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 570.00,898.50 A 28.50,28.50 0 0 1 541.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,870.00 A 28.50,28.50 0 0 1 630.00,841.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,870.00 A 28.50,28.50 0 0 1 630.00,898.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,870.00 A 28.50,28.50 0 0 1 690.00,841.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,870.00 A 28.50,28.50 0 0 1 690.00,898.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,898.50 A 28.50,28.50 0 0 1 721.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,841.50 A 28.50,28.50 0 0 1 778.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,870.00 A 28.50,28.50 0 0 1 810.00,898.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,870.00 A 28.50,28.50 0 0 1 810.00,841.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,841.50 A 28.50,28.50 0 0 1 898.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,898.50 A 28.50,28.50 0 0 1 841.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="870.0" fill="black" r="3.5999999999999996" /><path d="M 930.00,841.50 A 28.50,28.50 0 0 1 958.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,898.50 A 28.50,28.50 0 0 1 901.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,898.50 A 28.50,28.50 0 0 1 961.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,841.50 A 28.50,28.50 0 0 1 1018.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1050.00,841.50 A 28.50,28.50 0 0 1 1078.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1050.00,898.50 A 28.50,28.50 0 0 1 1021.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1050.0" cy="870.0" fill="black" r="3.5999999999999996" /><path d="M 1081.50,870.00 A 28.50,28.50 0 0 1 1110.00,841.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1138.50,870.00 A 28.50,28.50 0 0 1 1110.00,898.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1110.0" cy="870.0" fill="black" r="3.5999999999999996" /><path d="M 1141.50,870.00 A 28.50,28.50 0 0 1 1170.00,841.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,870.00 A 28.50,28.50 0 0 1 1170.00,898.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,898.50 A 28.50,28.50 0 0 1 1201.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,841.50 A 28.50,28.50 0 0 1 1258.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,870.00 A 28.50,28.50 0 0 1 1290.00,898.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,870.00 A 28.50,28.50 0 0 1 1290.00,841.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,841.50 A 28.50,28.50 0 0 1 1378.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,898.50 A 28.50,28.50 0 0 1 1321.50,870.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1350.0" cy="870.0" fill="black" r="3.5999999999999996" /><path d="M 150.00,901.50 A 28.50,28.50 0 0 1 178.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,958.50 A 28.50,28.50 0 0 1 121.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 238.50,930.00 A 28.50,28.50 0 0 1 210.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,930.00 A 28.50,28.50 0 0 1 210.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,958.50 A 28.50,28.50 0 0 1 241.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,901.50 A 28.50,28.50 0 0 1 298.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,958.50 A 28.50,28.50 0 0 1 301.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,901.50 A 28.50,28.50 0 0 1 358.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="330.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 361.50,930.00 A 28.50,28.50 0 0 1 390.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,930.00 A 28.50,28.50 0 0 1 390.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,930.00 A 28.50,28.50 0 0 1 450.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,930.00 A 28.50,28.50 0 0 1 450.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,901.50 A 28.50,28.50 0 0 1 538.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,958.50 A 28.50,28.50 0 0 1 481.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="510.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 541.50,930.00 A 28.50,28.50 0 0 1 570.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,930.00 A 28.50,28.50 0 0 1 570.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="570.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 601.50,930.00 A 28.50,28.50 0 0 1 630.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,930.00 A 28.50,28.50 0 0 1 630.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="630.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 661.50,930.00 A 28.50,28.50 0 0 1 690.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,930.00 A 28.50,28.50 0 0 1 690.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,901.50 A 28.50,28.50 0 0 1 778.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,958.50 A 28.50,28.50 0 0 1 721.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,930.00 A 28.50,28.50 0 0 1 810.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,930.00 A 28.50,28.50 0 0 1 810.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,930.00 A 28.50,28.50 0 0 1 870.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,930.00 A 28.50,28.50 0 0 1 870.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 958.50,930.00 A 28.50,28.50 0 0 1 930.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,930.00 A 28.50,28.50 0 0 1 930.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 990.00,901.50 A 28.50,28.50 0 0 1 1018.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,958.50 A 28.50,28.50 0 0 1 961.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="990.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 1021.50,930.00 A 28.50,28.50 0 0 1 1050.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,930.00 A 28.50,28.50 0 0 1 1050.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1050.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 1138.50,930.00 A 28.50,28.50 0 0 1 1110.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,930.00 A 28.50,28.50 0 0 1 1110.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,958.50 A 28.50,28.50 0 0 1 1141.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1170.00,901.50 A 28.50,28.50 0 0 1 1198.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,958.50 A 28.50,28.50 0 0 1 1201.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,901.50 A 28.50,28.50 0 0 1 1258.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1230.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 1290.00,901.50 A 28.50,28.50 0 0 1 1318.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,958.50 A 28.50,28.50 0 0 1 1261.50,930.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1290.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 1378.50,930.00 A 28.50,28.50 0 0 1 1350.00,958.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,930.00 A 28.50,28.50 0 0 1 1350.00,901.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1350.0" cy="930.0" fill="black" r="3.5999999999999996" /><path d="M 178.50,990.00 A 28.50,28.50 0 0 1 150.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 121.50,990.00 A 28.50,28.50 0 0 1 150.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 238.50,990.00 A 28.50,28.50 0 0 1 210.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,990.00 A 28.50,28.50 0 0 1 210.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="210.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 270.00,961.50 A 28.50,28.50 0 0 1 298.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,1018.50 A 28.50,28.50 0 0 1 241.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="270.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 301.50,990.00 A 28.50,28.50 0 0 1 330.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,990.00 A 28.50,28.50 0 0 1 330.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="330.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 418.50,990.00 A 28.50,28.50 0 0 1 390.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,990.00 A 28.50,28.50 0 0 1 390.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,1018.50 A 28.50,28.50 0 0 1 421.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 450.00,961.50 A 28.50,28.50 0 0 1 478.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,961.50 A 28.50,28.50 0 0 1 538.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 510.00,1018.50 A 28.50,28.50 0 0 1 481.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,990.00 A 28.50,28.50 0 0 1 570.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,990.00 A 28.50,28.50 0 0 1 570.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="570.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 630.00,1018.50 A 28.50,28.50 0 0 1 601.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,961.50 A 28.50,28.50 0 0 1 658.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,1018.50 A 28.50,28.50 0 0 1 661.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 690.00,961.50 A 28.50,28.50 0 0 1 718.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="690.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 750.00,961.50 A 28.50,28.50 0 0 1 778.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 750.00,1018.50 A 28.50,28.50 0 0 1 721.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="750.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 838.50,990.00 A 28.50,28.50 0 0 1 810.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,990.00 A 28.50,28.50 0 0 1 810.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,990.00 A 28.50,28.50 0 0 1 870.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,990.00 A 28.50,28.50 0 0 1 870.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,1018.50 A 28.50,28.50 0 0 1 901.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 930.00,961.50 A 28.50,28.50 0 0 1 958.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,961.50 A 28.50,28.50 0 0 1 1018.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,1018.50 A 28.50,28.50 0 0 1 961.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="990.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 1021.50,990.00 A 28.50,28.50 0 0 1 1050.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,990.00 A 28.50,28.50 0 0 1 1050.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1050.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 1138.50,990.00 A 28.50,28.50 0 0 1 1110.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,990.00 A 28.50,28.50 0 0 1 1110.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,990.00 A 28.50,28.50 0 0 1 1170.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1141.50,990.00 A 28.50,28.50 0 0 1 1170.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1170.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 1230.00,961.50 A 28.50,28.50 0 0 1 1258.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1230.00,1018.50 A 28.50,28.50 0 0 1 1201.50,990.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1230.0" cy="990.0" fill="black" r="3.5999999999999996" /><path d="M 1318.50,990.00 A 28.50,28.50 0 0 1 1290.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,990.00 A 28.50,28.50 0 0 1 1290.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,990.00 A 28.50,28.50 0 0 1 1350.00,1018.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,990.00 A 28.50,28.50 0 0 1 1350.00,961.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,1078.50 A 28.50,28.50 0 0 1 121.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,1021.50 A 28.50,28.50 0 0 1 178.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 210.00,1021.50 A 28.50,28.50 0 0 1 238.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 210.00,1078.50 A 28.50,28.50 0 0 1 181.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="210.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 241.50,1050.00 A 28.50,28.50 0 0 1 270.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 298.50,1050.00 A 28.50,28.50 0 0 1 270.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="270.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 330.00,1078.50 A 28.50,28.50 0 0 1 301.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,1021.50 A 28.50,28.50 0 0 1 358.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,1021.50 A 28.50,28.50 0 0 1 418.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 390.00,1078.50 A 28.50,28.50 0 0 1 361.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,1050.00 A 28.50,28.50 0 0 1 450.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,1050.00 A 28.50,28.50 0 0 1 450.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="450.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 481.50,1050.00 A 28.50,28.50 0 0 1 510.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 538.50,1050.00 A 28.50,28.50 0 0 1 510.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,1050.00 A 28.50,28.50 0 0 1 570.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,1050.00 A 28.50,28.50 0 0 1 570.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,1078.50 A 28.50,28.50 0 0 1 601.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,1021.50 A 28.50,28.50 0 0 1 658.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,1050.00 A 28.50,28.50 0 0 1 690.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,1050.00 A 28.50,28.50 0 0 1 690.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="690.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 721.50,1050.00 A 28.50,28.50 0 0 1 750.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 778.50,1050.00 A 28.50,28.50 0 0 1 750.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="750.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 838.50,1050.00 A 28.50,28.50 0 0 1 810.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,1050.00 A 28.50,28.50 0 0 1 810.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,1021.50 A 28.50,28.50 0 0 1 898.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,1078.50 A 28.50,28.50 0 0 1 841.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,1050.00 A 28.50,28.50 0 0 1 930.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,1050.00 A 28.50,28.50 0 0 1 930.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="930.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 961.50,1050.00 A 28.50,28.50 0 0 1 990.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1018.50,1050.00 A 28.50,28.50 0 0 1 990.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,1050.00 A 28.50,28.50 0 0 1 1050.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,1050.00 A 28.50,28.50 0 0 1 1050.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,1078.50 A 28.50,28.50 0 0 1 1081.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,1021.50 A 28.50,28.50 0 0 1 1138.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1110.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 1141.50,1050.00 A 28.50,28.50 0 0 1 1170.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,1050.00 A 28.50,28.50 0 0 1 1170.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1170.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 1201.50,1050.00 A 28.50,28.50 0 0 1 1230.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,1050.00 A 28.50,28.50 0 0 1 1230.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1230.0" cy="1050.0" fill="black" r="3.5999999999999996" /><path d="M 1290.00,1078.50 A 28.50,28.50 0 0 1 1261.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,1021.50 A 28.50,28.50 0 0 1 1318.50,1050.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,1050.00 A 28.50,28.50 0 0 1 1350.00,1078.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,1050.00 A 28.50,28.50 0 0 1 1350.00,1021.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,1081.50 A 28.50,28.50 0 0 1 178.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 150.00,1138.50 A 28.50,28.50 0 0 1 121.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="150.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 181.50,1110.00 A 28.50,28.50 0 0 1 210.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 238.50,1110.00 A 28.50,28.50 0 0 1 210.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="210.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 270.00,1138.50 A 28.50,28.50 0 0 1 241.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 270.00,1081.50 A 28.50,28.50 0 0 1 298.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,1138.50 A 28.50,28.50 0 0 1 301.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 330.00,1081.50 A 28.50,28.50 0 0 1 358.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,1110.00 A 28.50,28.50 0 0 1 390.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,1110.00 A 28.50,28.50 0 0 1 390.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="390.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 421.50,1110.00 A 28.50,28.50 0 0 1 450.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,1110.00 A 28.50,28.50 0 0 1 450.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 538.50,1110.00 A 28.50,28.50 0 0 1 510.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 481.50,1110.00 A 28.50,28.50 0 0 1 510.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,1110.00 A 28.50,28.50 0 0 1 570.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,1110.00 A 28.50,28.50 0 0 1 570.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,1081.50 A 28.50,28.50 0 0 1 658.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 630.00,1138.50 A 28.50,28.50 0 0 1 601.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="630.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 718.50,1110.00 A 28.50,28.50 0 0 1 690.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,1110.00 A 28.50,28.50 0 0 1 690.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 778.50,1110.00 A 28.50,28.50 0 0 1 750.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,1110.00 A 28.50,28.50 0 0 1 750.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,1110.00 A 28.50,28.50 0 0 1 810.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,1110.00 A 28.50,28.50 0 0 1 810.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="810.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 870.00,1081.50 A 28.50,28.50 0 0 1 898.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 870.00,1138.50 A 28.50,28.50 0 0 1 841.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="870.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 958.50,1110.00 A 28.50,28.50 0 0 1 930.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,1110.00 A 28.50,28.50 0 0 1 930.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,1081.50 A 28.50,28.50 0 0 1 1018.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 990.00,1138.50 A 28.50,28.50 0 0 1 961.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="990.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 1078.50,1110.00 A 28.50,28.50 0 0 1 1050.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,1110.00 A 28.50,28.50 0 0 1 1050.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1050.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 1110.00,1081.50 A 28.50,28.50 0 0 1 1138.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1110.00,1138.50 A 28.50,28.50 0 0 1 1081.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,1110.00 A 28.50,28.50 0 0 1 1170.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1141.50,1110.00 A 28.50,28.50 0 0 1 1170.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,1110.00 A 28.50,28.50 0 0 1 1230.00,1138.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1201.50,1110.00 A 28.50,28.50 0 0 1 1230.00,1081.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1230.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 1290.00,1138.50 A 28.50,28.50 0 0 1 1261.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1290.00,1081.50 A 28.50,28.50 0 0 1 1318.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1290.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 1350.00,1138.50 A 28.50,28.50 0 0 1 1321.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1350.00,1081.50 A 28.50,28.50 0 0 1 1378.50,1110.00" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><circle cx="1350.0" cy="1110.0" fill="black" r="3.5999999999999996" /><path d="M 178.50,1170.00 A 28.50,28.50 0 0 1 150.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 121.50,1170.00 A 28.50,28.50 0 0 1 150.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,1170.00 A 28.50,28.50 0 0 1 210.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 238.50,1170.00 A 28.50,28.50 0 0 1 210.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 241.50,1170.00 A 28.50,28.50 0 0 1 270.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 298.50,1170.00 A 28.50,28.50 0 0 1 270.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,1170.00 A 28.50,28.50 0 0 1 330.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,1170.00 A 28.50,28.50 0 0 1 330.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,1170.00 A 28.50,28.50 0 0 1 390.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,1170.00 A 28.50,28.50 0 0 1 390.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,1170.00 A 28.50,28.50 0 0 1 450.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,1170.00 A 28.50,28.50 0 0 1 450.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 481.50,1170.00 A 28.50,28.50 0 0 1 510.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 538.50,1170.00 A 28.50,28.50 0 0 1 510.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,1170.00 A 28.50,28.50 0 0 1 570.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,1170.00 A 28.50,28.50 0 0 1 570.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,1170.00 A 28.50,28.50 0 0 1 630.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,1170.00 A 28.50,28.50 0 0 1 630.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,1170.00 A 28.50,28.50 0 0 1 690.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,1170.00 A 28.50,28.50 0 0 1 690.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,1170.00 A 28.50,28.50 0 0 1 750.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 778.50,1170.00 A 28.50,28.50 0 0 1 750.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,1170.00 A 28.50,28.50 0 0 1 810.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,1170.00 A 28.50,28.50 0 0 1 810.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,1170.00 A 28.50,28.50 0 0 1 870.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,1170.00 A 28.50,28.50 0 0 1 870.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,1170.00 A 28.50,28.50 0 0 1 930.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,1170.00 A 28.50,28.50 0 0 1 930.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 961.50,1170.00 A 28.50,28.50 0 0 1 990.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1018.50,1170.00 A 28.50,28.50 0 0 1 990.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,1170.00 A 28.50,28.50 0 0 1 1050.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,1170.00 A 28.50,28.50 0 0 1 1050.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,1170.00 A 28.50,28.50 0 0 1 1110.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1138.50,1170.00 A 28.50,28.50 0 0 1 1110.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1141.50,1170.00 A 28.50,28.50 0 0 1 1170.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,1170.00 A 28.50,28.50 0 0 1 1170.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1201.50,1170.00 A 28.50,28.50 0 0 1 1230.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,1170.00 A 28.50,28.50 0 0 1 1230.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,1170.00 A 28.50,28.50 0 0 1 1290.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,1170.00 A 28.50,28.50 0 0 1 1290.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,1170.00 A 28.50,28.50 0 0 1 1350.00,1141.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,1170.00 A 28.50,28.50 0 0 1 1350.00,1198.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 121.50,1230.00 A 28.50,28.50 0 0 1 150.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 178.50,1230.00 A 28.50,28.50 0 0 1 150.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,1230.00 A 28.50,28.50 0 0 1 210.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 238.50,1230.00 A 28.50,28.50 0 0 1 210.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 241.50,1230.00 A 28.50,28.50 0 0 1 270.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 298.50,1230.00 A 28.50,28.50 0 0 1 270.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,1230.00 A 28.50,28.50 0 0 1 330.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,1230.00 A 28.50,28.50 0 0 1 330.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,1230.00 A 28.50,28.50 0 0 1 390.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,1230.00 A 28.50,28.50 0 0 1 390.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,1230.00 A 28.50,28.50 0 0 1 450.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,1230.00 A 28.50,28.50 0 0 1 450.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 481.50,1230.00 A 28.50,28.50 0 0 1 510.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 538.50,1230.00 A 28.50,28.50 0 0 1 510.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,1230.00 A 28.50,28.50 0 0 1 570.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,1230.00 A 28.50,28.50 0 0 1 570.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,1230.00 A 28.50,28.50 0 0 1 630.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,1230.00 A 28.50,28.50 0 0 1 630.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,1230.00 A 28.50,28.50 0 0 1 690.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,1230.00 A 28.50,28.50 0 0 1 690.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,1230.00 A 28.50,28.50 0 0 1 750.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 778.50,1230.00 A 28.50,28.50 0 0 1 750.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,1230.00 A 28.50,28.50 0 0 1 810.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,1230.00 A 28.50,28.50 0 0 1 810.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,1230.00 A 28.50,28.50 0 0 1 870.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,1230.00 A 28.50,28.50 0 0 1 870.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,1230.00 A 28.50,28.50 0 0 1 930.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,1230.00 A 28.50,28.50 0 0 1 930.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 961.50,1230.00 A 28.50,28.50 0 0 1 990.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1018.50,1230.00 A 28.50,28.50 0 0 1 990.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,1230.00 A 28.50,28.50 0 0 1 1050.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,1230.00 A 28.50,28.50 0 0 1 1050.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,1230.00 A 28.50,28.50 0 0 1 1110.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1138.50,1230.00 A 28.50,28.50 0 0 1 1110.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1141.50,1230.00 A 28.50,28.50 0 0 1 1170.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,1230.00 A 28.50,28.50 0 0 1 1170.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1201.50,1230.00 A 28.50,28.50 0 0 1 1230.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,1230.00 A 28.50,28.50 0 0 1 1230.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,1230.00 A 28.50,28.50 0 0 1 1290.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,1230.00 A 28.50,28.50 0 0 1 1290.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,1230.00 A 28.50,28.50 0 0 1 1350.00,1201.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,1230.00 A 28.50,28.50 0 0 1 1350.00,1258.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 121.50,1290.00 A 28.50,28.50 0 0 1 150.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 178.50,1290.00 A 28.50,28.50 0 0 1 150.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,1290.00 A 28.50,28.50 0 0 1 210.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 238.50,1290.00 A 28.50,28.50 0 0 1 210.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 241.50,1290.00 A 28.50,28.50 0 0 1 270.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 298.50,1290.00 A 28.50,28.50 0 0 1 270.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,1290.00 A 28.50,28.50 0 0 1 330.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,1290.00 A 28.50,28.50 0 0 1 330.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,1290.00 A 28.50,28.50 0 0 1 390.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,1290.00 A 28.50,28.50 0 0 1 390.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,1290.00 A 28.50,28.50 0 0 1 450.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,1290.00 A 28.50,28.50 0 0 1 450.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 481.50,1290.00 A 28.50,28.50 0 0 1 510.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 538.50,1290.00 A 28.50,28.50 0 0 1 510.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,1290.00 A 28.50,28.50 0 0 1 570.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,1290.00 A 28.50,28.50 0 0 1 570.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,1290.00 A 28.50,28.50 0 0 1 630.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,1290.00 A 28.50,28.50 0 0 1 630.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,1290.00 A 28.50,28.50 0 0 1 690.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,1290.00 A 28.50,28.50 0 0 1 690.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,1290.00 A 28.50,28.50 0 0 1 750.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 778.50,1290.00 A 28.50,28.50 0 0 1 750.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,1290.00 A 28.50,28.50 0 0 1 810.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,1290.00 A 28.50,28.50 0 0 1 810.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,1290.00 A 28.50,28.50 0 0 1 870.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,1290.00 A 28.50,28.50 0 0 1 870.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,1290.00 A 28.50,28.50 0 0 1 930.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,1290.00 A 28.50,28.50 0 0 1 930.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 961.50,1290.00 A 28.50,28.50 0 0 1 990.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1018.50,1290.00 A 28.50,28.50 0 0 1 990.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,1290.00 A 28.50,28.50 0 0 1 1050.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,1290.00 A 28.50,28.50 0 0 1 1050.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,1290.00 A 28.50,28.50 0 0 1 1110.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1138.50,1290.00 A 28.50,28.50 0 0 1 1110.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1141.50,1290.00 A 28.50,28.50 0 0 1 1170.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,1290.00 A 28.50,28.50 0 0 1 1170.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1201.50,1290.00 A 28.50,28.50 0 0 1 1230.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,1290.00 A 28.50,28.50 0 0 1 1230.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,1290.00 A 28.50,28.50 0 0 1 1290.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,1290.00 A 28.50,28.50 0 0 1 1290.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,1290.00 A 28.50,28.50 0 0 1 1350.00,1261.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,1290.00 A 28.50,28.50 0 0 1 1350.00,1318.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 121.50,1350.00 A 28.50,28.50 0 0 1 150.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 178.50,1350.00 A 28.50,28.50 0 0 1 150.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 181.50,1350.00 A 28.50,28.50 0 0 1 210.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 238.50,1350.00 A 28.50,28.50 0 0 1 210.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 241.50,1350.00 A 28.50,28.50 0 0 1 270.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 298.50,1350.00 A 28.50,28.50 0 0 1 270.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 301.50,1350.00 A 28.50,28.50 0 0 1 330.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 358.50,1350.00 A 28.50,28.50 0 0 1 330.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 361.50,1350.00 A 28.50,28.50 0 0 1 390.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 418.50,1350.00 A 28.50,28.50 0 0 1 390.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 421.50,1350.00 A 28.50,28.50 0 0 1 450.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 478.50,1350.00 A 28.50,28.50 0 0 1 450.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 481.50,1350.00 A 28.50,28.50 0 0 1 510.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 538.50,1350.00 A 28.50,28.50 0 0 1 510.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 541.50,1350.00 A 28.50,28.50 0 0 1 570.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 598.50,1350.00 A 28.50,28.50 0 0 1 570.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 601.50,1350.00 A 28.50,28.50 0 0 1 630.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 658.50,1350.00 A 28.50,28.50 0 0 1 630.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 661.50,1350.00 A 28.50,28.50 0 0 1 690.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 718.50,1350.00 A 28.50,28.50 0 0 1 690.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 721.50,1350.00 A 28.50,28.50 0 0 1 750.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 778.50,1350.00 A 28.50,28.50 0 0 1 750.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 781.50,1350.00 A 28.50,28.50 0 0 1 810.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 838.50,1350.00 A 28.50,28.50 0 0 1 810.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 841.50,1350.00 A 28.50,28.50 0 0 1 870.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 898.50,1350.00 A 28.50,28.50 0 0 1 870.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 901.50,1350.00 A 28.50,28.50 0 0 1 930.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 958.50,1350.00 A 28.50,28.50 0 0 1 930.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 961.50,1350.00 A 28.50,28.50 0 0 1 990.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1018.50,1350.00 A 28.50,28.50 0 0 1 990.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1021.50,1350.00 A 28.50,28.50 0 0 1 1050.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1078.50,1350.00 A 28.50,28.50 0 0 1 1050.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1081.50,1350.00 A 28.50,28.50 0 0 1 1110.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1138.50,1350.00 A 28.50,28.50 0 0 1 1110.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1141.50,1350.00 A 28.50,28.50 0 0 1 1170.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1198.50,1350.00 A 28.50,28.50 0 0 1 1170.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1201.50,1350.00 A 28.50,28.50 0 0 1 1230.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1258.50,1350.00 A 28.50,28.50 0 0 1 1230.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1261.50,1350.00 A 28.50,28.50 0 0 1 1290.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1318.50,1350.00 A 28.50,28.50 0 0 1 1290.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1321.50,1350.00 A 28.50,28.50 0 0 1 1350.00,1321.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /><path d="M 1378.50,1350.00 A 28.50,28.50 0 0 1 1350.00,1378.50" fill="none" stroke="black" stroke-linecap="round" stroke-width="1.7" /></g></svg>